package constelation is

  constant constelationName : string := "IRNSSL5";

  constant radioFrequencyOut : integer := 1176450000;
  constant outputRate        : integer := 1023000;--2600000;

  constant RadioFrequencyIn : integer := 1176450000;
  constant InputRate        : integer := 1023000;
  constant FrameSize        : integer := 5;

end package;