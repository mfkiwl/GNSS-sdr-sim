library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package input is
  
  constant inputFrameSatCount : integer := 1;
  
  type inputTable is array(0 to 100 - 1) of std_logic_vector(176-1 downto 0);
  constant inputSeq : inputTable := (
    x"000600000000000000070000000000000000000000ff",
    x"000600000000000000120000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000140000000000000000000000ff",
    x"0006000000000000000a0000000000000000000000ff",
    x"000600000000000000090000000000000000000000ff",
    x"000600000000000000040000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000180000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000100000000000000000000000ff",
    x"000600000000000000130000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"0006000000000000000a0000000000000000000000ff",
    x"000600000000000000110000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"000600000000000000180000000000000000000000ff",
    x"000600000000000000100000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"000600000000000000110000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000150000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"000600000000000000050000000000000000000000ff",
    x"000600000000000000050000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000010000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000040000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000010000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000140000000000000000000000ff",
    x"000600000000000000180000000000000000000000ff",
    x"0006000000000000001e0000000000000000000000ff",
    x"000600000000000000070000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"000600000000000000190000000000000000000000ff",
    x"000600000000000000070000000000000000000000ff",
    x"0006000000000000001a0000000000000000000000ff",
    x"000600000000000000130000000000000000000000ff",
    x"000600000000000000170000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000120000000000000000000000ff",
    x"000600000000000000190000000000000000000000ff",
    x"000600000000000000070000000000000000000000ff",
    x"000600000000000000120000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000120000000000000000000000ff",
    x"0006000000000000000a0000000000000000000000ff",
    x"000600000000000000010000000000000000000000ff",
    x"000600000000000000040000000000000000000000ff",
    x"000600000000000000000000000000000000000000ff",
    x"000600000000000000120000000000000000000000ff",
    x"000600000000000000190000000000000000000000ff",
    x"000600000000000000030000000000000000000000ff",
    x"0006000000000000000b0000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"000600000000000000100000000000000000000000ff",
    x"000600000000000000010000000000000000000000ff",
    x"000600000000000000010000000000000000000000ff",
    x"000600000000000000040000000000000000000000ff",
    x"000600000000000000130000000000000000000000ff",
    x"0006000000000000001c0000000000000000000000ff",
    x"000600000000000000020000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000150000000000000000000000ff",
    x"0006000000000000001d0000000000000000000000ff",
    x"0006000000000000001a0000000000000000000000ff",
    x"000600000000000000070000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000110000000000000000000000ff",
    x"000600000000000000140000000000000000000000ff",
    x"000600000000000000030000000000000000000000ff",
    x"000600000000000000080000000000000000000000ff",
    x"000600000000000000170000000000000000000000ff",
    x"000600000000000000030000000000000000000000ff",
    x"000600000000000000150000000000000000000000ff",
    x"0006000000000000000b0000000000000000000000ff",
    x"0006000000000000000c0000000000000000000000ff",
    x"0006000000000000001b0000000000000000000000ff",
    x"000600000000000000120000000000000000000000ff",
    x"000600000000000000180000000000000000000000ff",
    x"0006000000000000000c0000000000000000000000ff",
    x"000600000000000000170000000000000000000000ff"
  );
end package;