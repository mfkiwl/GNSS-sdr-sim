library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package input is
  
  constant inputFrameSatCount : integer := 25;
  
  type inputTable is array(0 to 50424 - 1) of std_logic_vector(176-1 downto 0);
  constant inputSeq : inputTable := (
    x"000100000000000001aa000000002f57460266e3681c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa000000003c8d8a0bfbe5401c",
    x"020900000000000001aa00000000396528fb33889b1c",
    x"030b00000000000001aa000000003d37110003e39f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aa0000000035d394099dd2cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa00000000331c7f072f4bc51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa000000002f31b404cd3c411c",
    x"070a00000000000001aa0000000039a909ef36078a1c",
    x"080200000000000001aa00000000360aeaf669ec871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266e3641c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe5411c",
    x"0209000000000000029500000000000000fb3388951c",
    x"030b0000000000000295fffffffffffff50003e3a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd2c91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4bc21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd3c3b1c",
    x"070a0000000000000295fffffffffffff8ef3607871c",
    x"08020000000000000295fffffffffffff6f669ec841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266e3601c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe5421c",
    x"0209000000000000015a00000000000000fb33888f1c",
    x"030b000000000000015afffffffffffff50003e3a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dd2c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f4bbe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd3c351c",
    x"070a000000000000015afffffffffffff8ef3607831c",
    x"0802000000000000015afffffffffffff6f669ec821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e35b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5431c",
    x"0209000000000000015500000000000000fb33888a1c",
    x"030b0000000000000155fffffffffffff50003e3a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd2c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4bba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3c2f1c",
    x"070a0000000000000155fffffffffffff8ef3607801c",
    x"08020000000000000155fffffffffffff6f669ec801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266e3571c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe5441c",
    x"020900000000000002a900000000000000fb3388841c",
    x"030b0000000000000155fffffffffffff50003e3a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd2c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4bb61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd3c291c",
    x"070a0000000000000155fffffffffffff8ef36077c1c",
    x"080200000000000002a9fffffffffffff6f669ec7d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266e3531c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5461c",
    x"0209000000000000029a00000000000000fb33887f1c",
    x"030b0000000000000265fffffffffffff50003e3a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dd2c01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f4bb31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd3c231c",
    x"070a0000000000000255fffffffffffff8ef3607781c",
    x"080200000000000002a9fffffffffffff6f669ec7b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e34f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe5471c",
    x"0209000000000000015a00000000000000fb3388791c",
    x"030b0000000000000265fffffffffffff50003e3a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dd2be1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4baf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd3c1d1c",
    x"070a000000000000029afffffffffffff8ef3607751c",
    x"0802000000000000019afffffffffffff6f669ec791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266e34b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe5481c",
    x"0209000000000000019900000000000000fb3388731c",
    x"030b0000000000000166fffffffffffff50003e3a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dd2bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f4bab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd3c161c",
    x"070a00000000000001a9fffffffffffff8ef3607711c",
    x"0802000000000000026afffffffffffff6f669ec761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266e3461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002690000000000000b0bfbe5491c",
    x"0209000000000000016600000000000000fb33886e1c",
    x"030b00000000000001a6fffffffffffff50003e3a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dd2b91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f4ba71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd3c101c",
    x"070a0000000000000199fffffffffffff8ef36076e1c",
    x"0802000000000000025afffffffffffff6f669ec741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266e3421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe54a1c",
    x"0209000000000000015500000000000000fb3388681c",
    x"030b000000000000015afffffffffffff50003e3a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dd2b71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f4ba41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd3c0a1c",
    x"070a000000000000016afffffffffffff8ef36076a1c",
    x"0802000000000000025afffffffffffff6f669ec721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266e33e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe54b1c",
    x"0209000000000000015a00000000000000fb3388631c",
    x"030b0000000000000295fffffffffffff50003e3a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2b41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f4ba01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd3c041c",
    x"070a00000000000001aafffffffffffff8ef3607671c",
    x"08020000000000000296fffffffffffff6f669ec6f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266e33a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002990000000000000b0bfbe54c1c",
    x"020900000000000001a900000000000000fb33885d1c",
    x"030b0000000000000299fffffffffffff50003e3ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dd2b21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f4b9c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd3bfe1c",
    x"070a0000000000000165fffffffffffff8ef3607631c",
    x"0802000000000000016afffffffffffff6f669ec6d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266e3361c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe54d1c",
    x"020900000000000002aa00000000000000fb3388581c",
    x"030b0000000000000169fffffffffffff50003e3ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dd2b01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd3bf81c",
    x"070a00000000000002a9fffffffffffff8ef3607601c",
    x"08020000000000000199fffffffffffff6f669ec6a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000299ffffffffffffff0266e3311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe54e1c",
    x"0209000000000000029a00000000000000fb3388521c",
    x"030b000000000000019afffffffffffff50003e3ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dd2ad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b951c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd3bf21c",
    x"070a000000000000016afffffffffffff8ef36075c1c",
    x"08020000000000000165fffffffffffff6f669ec681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266e32d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe54f1c",
    x"020900000000000002a600000000000000fb33884c1c",
    x"030b000000000000015afffffffffffff50003e3ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dd2ab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd3bec1c",
    x"070a000000000000025afffffffffffff8ef3607591c",
    x"0802000000000000025afffffffffffff6f669ec661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266e3291c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe5501c",
    x"0209000000000000015a00000000000000fb3388471c",
    x"030b0000000000000195fffffffffffff50003e3af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dd2a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002990000000000000b072f4b8d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026affffffffffffff04cd3be51c",
    x"070a00000000000002a9fffffffffffff8ef3607551c",
    x"08020000000000000259fffffffffffff6f669ec631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266e3251c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe5511c",
    x"020900000000000002a600000000000000fb3388411c",
    x"030b0000000000000159fffffffffffff50003e3b01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dd2a61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4b891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd3bdf1c",
    x"070a0000000000000159fffffffffffff8ef3607521c",
    x"08020000000000000295fffffffffffff6f669ec611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e3211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5531c",
    x"0209000000000000031f00000000000000fb33883c1c",
    x"030b000000000000031ffffffffffffff50003e3b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd2a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f4b861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd3bd91c",
    x"070a000000000000031ffffffffffffff8ef36074e1c",
    x"0802000000000000031ffffffffffffff6f669ec5f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e31c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5541c",
    x"020900000000000000ae00000000000000fb3388361c",
    x"030b00000000000000aefffffffffffff50003e3b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd2a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f4b821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd3bd31c",
    x"070a00000000000000aefffffffffffff8ef36074a1c",
    x"080200000000000000aefffffffffffff6f669ec5c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e3181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5551c",
    x"020900000000000001a400000000000000fb3388301c",
    x"030b00000000000001a4fffffffffffff50003e3b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd29f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f4b7e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd3bcd1c",
    x"070a00000000000001a4fffffffffffff8ef3607471c",
    x"080200000000000001a4fffffffffffff6f669ec5a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e3141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe5561c",
    x"0209000000000000016a00000000000000fb33882b1c",
    x"030b000000000000016afffffffffffff50003e3b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dd29d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f4b7a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd3bc71c",
    x"070a000000000000016afffffffffffff8ef3607431c",
    x"0802000000000000016afffffffffffff6f669ec571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e3101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5571c",
    x"0209000000000000015500000000000000fb3388251c",
    x"030b0000000000000155fffffffffffff50003e3b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd29a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4b771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3bc11c",
    x"070a0000000000000155fffffffffffff8ef3607401c",
    x"08020000000000000155fffffffffffff6f669ec551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266e30b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe5581c",
    x"0209000000000000019500000000000000fb3388201c",
    x"030b0000000000000195fffffffffffff50003e3b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dd2981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f4b731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd3bbb1c",
    x"070a0000000000000195fffffffffffff8ef36073c1c",
    x"080200000000000002a5fffffffffffff6f669ec531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e3071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5591c",
    x"020900000000000002aa00000000000000fb33881a1c",
    x"030b00000000000002aafffffffffffff50003e3b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4b6f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3bb41c",
    x"070a00000000000002aafffffffffffff8ef3607391c",
    x"08020000000000000155fffffffffffff6f669ec501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266e3031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe55a1c",
    x"0209000000000000029600000000000000fb3388141c",
    x"030b00000000000001aafffffffffffff50003e3b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dd2931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4b6c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd3bae1c",
    x"070a0000000000000256fffffffffffff8ef3607351c",
    x"08020000000000000155fffffffffffff6f669ec4e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266e2ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe55b1c",
    x"0209000000000000026500000000000000fb33880f1c",
    x"030b00000000000002a9fffffffffffff50003e3b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dd2911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f4b681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd3ba81c",
    x"070a000000000000029afffffffffffff8ef3607321c",
    x"08020000000000000159fffffffffffff6f669ec4c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266e2fb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe55c1c",
    x"0209000000000000029600000000000000fb3388091c",
    x"030b000000000000016afffffffffffff50003e3ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dd28f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f4b641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd3ba21c",
    x"070a0000000000000159fffffffffffff8ef36072e1c",
    x"0802000000000000015afffffffffffff6f669ec491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266e2f61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe55d1c",
    x"0209000000000000016900000000000000fb3388041c",
    x"030b0000000000000295fffffffffffff50003e3bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dd28c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b601c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd3b9c1c",
    x"070a0000000000000196fffffffffffff8ef36072b1c",
    x"08020000000000000299fffffffffffff6f669ec471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e2f21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe55e1c",
    x"020900000000000002a500000000000000fb3387fe1c",
    x"030b0000000000000156fffffffffffff50003e3bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dd28a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f4b5d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd3b961c",
    x"070a00000000000002a6fffffffffffff8ef3607271c",
    x"080200000000000001a5fffffffffffff6f669ec451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266e2ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe5601c",
    x"0209000000000000025500000000000000fb3387f91c",
    x"030b000000000000016afffffffffffff50003e3be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dd2881c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f4b591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd3b901c",
    x"070a0000000000000295fffffffffffff8ef3607231c",
    x"0802000000000000026afffffffffffff6f669ec421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266e2ea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe5611c",
    x"0209000000000000029a00000000000000fb3387f31c",
    x"030b0000000000000269fffffffffffff50003e3bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dd2851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f4b551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd3b8a1c",
    x"070a0000000000000196fffffffffffff8ef3607201c",
    x"08020000000000000165fffffffffffff6f669ec401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2e61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe5621c",
    x"020900000000000001a600000000000000fb3387ed1c",
    x"030b000000000000019afffffffffffff50003e3c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dd2831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f4b511c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd3b831c",
    x"070a000000000000026afffffffffffff8ef36071c1c",
    x"0802000000000000019afffffffffffff6f669ec3d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266e2e11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbe5631c",
    x"0209000000000000025a00000000000000fb3387e81c",
    x"030b00000000000002a9fffffffffffff50003e3c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dd2811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f4b4e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd3b7d1c",
    x"070a00000000000002a6fffffffffffff8ef3607191c",
    x"08020000000000000295fffffffffffff6f669ec3b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266e2dd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe5641c",
    x"0209000000000000029600000000000000fb3387e21c",
    x"030b000000000000025afffffffffffff50003e3c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dd27e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f4b4a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd3b771c",
    x"070a000000000000019afffffffffffff8ef3607151c",
    x"0802000000000000029afffffffffffff6f669ec391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266e2d91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe5651c",
    x"0209000000000000019900000000000000fb3387dd1c",
    x"030b0000000000000156fffffffffffff50003e3c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd27c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f4b461c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd3b711c",
    x"070a0000000000000166fffffffffffff8ef3607121c",
    x"080200000000000001a9fffffffffffff6f669ec361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e2d51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe5661c",
    x"0209000000000000015600000000000000fb3387d71c",
    x"030b0000000000000169fffffffffffff50003e3c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dd27a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f4b421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd3b6b1c",
    x"070a0000000000000159fffffffffffff8ef36070e1c",
    x"08020000000000000255fffffffffffff6f669ec341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266e2d11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5671c",
    x"0209000000000000029a00000000000000fb3387d11c",
    x"030b00000000000002a9fffffffffffff50003e3c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dd2771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4b3f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd3b651c",
    x"070a0000000000000159fffffffffffff8ef36070b1c",
    x"08020000000000000299fffffffffffff6f669ec321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e2cc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5681c",
    x"0209000000000000031f00000000000000fb3387cc1c",
    x"030b000000000000031ffffffffffffff50003e3c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd2751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f4b3b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd3b5f1c",
    x"070a000000000000031ffffffffffffff8ef3607071c",
    x"0802000000000000031ffffffffffffff6f669ec2f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e2c81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5691c",
    x"020900000000000000ae00000000000000fb3387c61c",
    x"030b00000000000000aefffffffffffff50003e3c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd2731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f4b371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd3b591c",
    x"070a00000000000000aefffffffffffff8ef3607041c",
    x"080200000000000000aefffffffffffff6f669ec2d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e2c41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe56a1c",
    x"020900000000000001a400000000000000fb3387c11c",
    x"030b00000000000001a4fffffffffffff50003e3c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd2701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f4b331c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd3b521c",
    x"070a00000000000001a4fffffffffffff8ef3607001c",
    x"080200000000000001a4fffffffffffff6f669ec2b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266e2c01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe56b1c",
    x"0209000000000000026a00000000000000fb3387bb1c",
    x"030b000000000000026afffffffffffff50003e3c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dd26e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f4b301c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026affffffffffffff04cd3b4c1c",
    x"070a000000000000026afffffffffffff8ef3606fc1c",
    x"0802000000000000026afffffffffffff6f669ec281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e2bc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe56d1c",
    x"0209000000000000015500000000000000fb3387b61c",
    x"030b0000000000000155fffffffffffff50003e3ca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd26c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f4b2c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd3b461c",
    x"070a00000000000002a9fffffffffffff8ef3606f91c",
    x"08020000000000000155fffffffffffff6f669ec261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e2b71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe56e1c",
    x"0209000000000000015500000000000000fb3387b01c",
    x"030b0000000000000155fffffffffffff50003e3cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd2691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4b281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3b401c",
    x"070a00000000000001aafffffffffffff8ef3606f51c",
    x"08020000000000000155fffffffffffff6f669ec231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266e2b31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe56f1c",
    x"0209000000000000015600000000000000fb3387aa1c",
    x"030b0000000000000155fffffffffffff50003e3cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dd2671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f4b241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd3b3a1c",
    x"070a00000000000002aafffffffffffff8ef3606f21c",
    x"08020000000000000155fffffffffffff6f669ec211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e2af1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe5701c",
    x"0209000000000000025500000000000000fb3387a51c",
    x"030b0000000000000195fffffffffffff50003e3cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd2651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f4b211c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd3b341c",
    x"070a000000000000026afffffffffffff8ef3606ee1c",
    x"08020000000000000195fffffffffffff6f669ec1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266e2ab1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe5711c",
    x"0209000000000000016500000000000000fb33879f1c",
    x"030b00000000000002a9fffffffffffff50003e3cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dd2621c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4b1d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000259ffffffffffffff04cd3b2e1c",
    x"070a0000000000000256fffffffffffff8ef3606eb1c",
    x"08020000000000000299fffffffffffff6f669ec1c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266e2a61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe5721c",
    x"0209000000000000019900000000000000fb33879a1c",
    x"030b0000000000000195fffffffffffff50003e3d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dd2601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd3b281c",
    x"070a0000000000000266fffffffffffff8ef3606e71c",
    x"080200000000000002a6fffffffffffff6f669ec1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266e2a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe5731c",
    x"0209000000000000016500000000000000fb3387941c",
    x"030b0000000000000166fffffffffffff50003e3d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dd25e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f4b151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd3b221c",
    x"070a0000000000000156fffffffffffff8ef3606e41c",
    x"0802000000000000025afffffffffffff6f669ec181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266e29e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe5741c",
    x"0209000000000000019500000000000000fb33878e1c",
    x"030b0000000000000265fffffffffffff50003e3d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dd25b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd3b1b1c",
    x"070a000000000000025afffffffffffff8ef3606e01c",
    x"0802000000000000016afffffffffffff6f669ec151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e29a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe5751c",
    x"0209000000000000026a00000000000000fb3387891c",
    x"030b00000000000002aafffffffffffff50003e3d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd2591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f4b0e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd3b151c",
    x"070a0000000000000195fffffffffffff8ef3606dd1c",
    x"08020000000000000195fffffffffffff6f669ec131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266e2961c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe5761c",
    x"0209000000000000025600000000000000fb3387831c",
    x"030b00000000000002a5fffffffffffff50003e3d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dd2571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f4b0a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd3b0f1c",
    x"070a00000000000002a5fffffffffffff8ef3606d91c",
    x"08020000000000000295fffffffffffff6f669ec101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266e2911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe5771c",
    x"020900000000000001a900000000000000fb33877e1c",
    x"030b0000000000000155fffffffffffff50003e3d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dd2541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f4b071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd3b091c",
    x"070a0000000000000256fffffffffffff8ef3606d61c",
    x"08020000000000000199fffffffffffff6f669ec0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266e28d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe5781c",
    x"0209000000000000029500000000000000fb3387781c",
    x"030b0000000000000299fffffffffffff50003e3d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f4b031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd3b031c",
    x"070a0000000000000266fffffffffffff8ef3606d21c",
    x"08020000000000000166fffffffffffff6f669ec0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266e2891c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe57a1c",
    x"0209000000000000016900000000000000fb3387731c",
    x"030b000000000000016afffffffffffff50003e3d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dd2501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f4aff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd3afd1c",
    x"070a0000000000000256fffffffffffff8ef3606ce1c",
    x"08020000000000000199fffffffffffff6f669ec091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266e2851c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe57b1c",
    x"0209000000000000026a00000000000000fb33876d1c",
    x"030b000000000000016afffffffffffff50003e3d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dd24d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f4afb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd3af71c",
    x"070a00000000000001a5fffffffffffff8ef3606cb1c",
    x"08020000000000000266fffffffffffff6f669ec071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266e2811c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe57c1c",
    x"020900000000000001a900000000000000fb3387671c",
    x"030b000000000000026afffffffffffff50003e3d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dd24b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f4af81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd3af01c",
    x"070a0000000000000166fffffffffffff8ef3606c71c",
    x"08020000000000000296fffffffffffff6f669ec051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266e27c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe57d1c",
    x"020900000000000002a600000000000000fb3387621c",
    x"030b000000000000015afffffffffffff50003e3da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dd2491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f4af41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd3aea1c",
    x"070a0000000000000295fffffffffffff8ef3606c41c",
    x"080200000000000002a5fffffffffffff6f669ec021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e2781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe57e1c",
    x"0209000000000000031f00000000000000fb33875c1c",
    x"030b000000000000031ffffffffffffff50003e3db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd2461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f4af01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd3ae41c",
    x"070a000000000000031ffffffffffffff8ef3606c01c",
    x"0802000000000000031ffffffffffffff6f669ec001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e2741c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe57f1c",
    x"020900000000000000ae00000000000000fb3387571c",
    x"030b00000000000000aefffffffffffff50003e3dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd2441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f4aec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd3ade1c",
    x"070a00000000000000aefffffffffffff8ef3606bd1c",
    x"080200000000000000aefffffffffffff6f669ebfe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e2701c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5801c",
    x"020900000000000001a400000000000000fb3387511c",
    x"030b00000000000001a4fffffffffffff50003e3dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd2421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f4ae91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd3ad81c",
    x"070a00000000000001a4fffffffffffff8ef3606b91c",
    x"080200000000000001a4fffffffffffff6f669ebfb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266e26c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe5811c",
    x"0209000000000000015a00000000000000fb33874b1c",
    x"030b000000000000015afffffffffffff50003e3de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dd23f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f4ae51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd3ad21c",
    x"070a000000000000015afffffffffffff8ef3606b61c",
    x"0802000000000000015afffffffffffff6f669ebf91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5821c",
    x"020900000000000001aa00000000000000fb3387461c",
    x"030b0000000000000255fffffffffffff50003e3df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd23d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4ae11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3acc1c",
    x"070a0000000000000155fffffffffffff8ef3606b21c",
    x"08020000000000000155fffffffffffff6f669ebf61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266e2631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe5831c",
    x"0209000000000000016900000000000000fb3387401c",
    x"030b0000000000000269fffffffffffff50003e3e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dd23a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f4add1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd3ac61c",
    x"070a00000000000002a6fffffffffffff8ef3606af1c",
    x"080200000000000001a5fffffffffffff6f669ebf41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266e25f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe5841c",
    x"020900000000000001a600000000000000fb33873b1c",
    x"030b0000000000000296fffffffffffff50003e3e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dd2381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f4ada1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd3abf1c",
    x"070a000000000000029afffffffffffff8ef3606ab1c",
    x"08020000000000000196fffffffffffff6f669ebf21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266e25b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe5861c",
    x"0209000000000000026900000000000000fb3387351c",
    x"030b0000000000000255fffffffffffff50003e3e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dd2361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f4ad61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000199ffffffffffffff04cd3ab91c",
    x"070a0000000000000265fffffffffffff8ef3606a71c",
    x"08020000000000000256fffffffffffff6f669ebef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2571c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe5871c",
    x"0209000000000000015600000000000000fb3387301c",
    x"030b0000000000000155fffffffffffff50003e3e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f4ad21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd3ab31c",
    x"070a00000000000002aafffffffffffff8ef3606a41c",
    x"08020000000000000155fffffffffffff6f669ebed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266e2521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbe5881c",
    x"0209000000000000025500000000000000fb33872a1c",
    x"030b0000000000000255fffffffffffff50003e3e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dd2311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f4ace1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd3aad1c",
    x"070a00000000000001aafffffffffffff8ef3606a01c",
    x"08020000000000000255fffffffffffff6f669ebeb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e24e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5891c",
    x"0209000000000000015500000000000000fb3387241c",
    x"030b0000000000000155fffffffffffff50003e3e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd22f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4acb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3aa71c",
    x"070a00000000000002aafffffffffffff8ef36069d1c",
    x"08020000000000000155fffffffffffff6f669ebe81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e24a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe58a1c",
    x"0209000000000000015500000000000000fb33871f1c",
    x"030b0000000000000155fffffffffffff50003e3e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd22c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4ac71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3aa11c",
    x"070a00000000000002aafffffffffffff8ef3606991c",
    x"08020000000000000155fffffffffffff6f669ebe61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe58b1c",
    x"0209000000000000015500000000000000fb3387191c",
    x"030b0000000000000155fffffffffffff50003e3e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd22a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4ac31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a9b1c",
    x"070a00000000000002aafffffffffffff8ef3606961c",
    x"08020000000000000155fffffffffffff6f669ebe31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266e2421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe58c1c",
    x"0209000000000000025900000000000000fb3387141c",
    x"030b0000000000000259fffffffffffff50003e3e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dd2281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f4ac01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000259ffffffffffffff04cd3a951c",
    x"070a00000000000001a6fffffffffffff8ef3606921c",
    x"08020000000000000259fffffffffffff6f669ebe11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e23d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe58d1c",
    x"0209000000000000015500000000000000fb33870e1c",
    x"030b0000000000000155fffffffffffff50003e3ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4abc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a8e1c",
    x"070a00000000000002aafffffffffffff8ef36068f1c",
    x"08020000000000000155fffffffffffff6f669ebdf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe58e1c",
    x"0209000000000000015500000000000000fb3387081c",
    x"030b0000000000000155fffffffffffff50003e3eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4ab81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a881c",
    x"070a00000000000002aafffffffffffff8ef36068b1c",
    x"08020000000000000155fffffffffffff6f669ebdc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266e2351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbe58f1c",
    x"0209000000000000015900000000000000fb3387031c",
    x"030b0000000000000159fffffffffffff50003e3ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dd2211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f4ab41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd3a821c",
    x"070a00000000000002a6fffffffffffff8ef3606871c",
    x"08020000000000000159fffffffffffff6f669ebda1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266e2311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe5901c",
    x"0209000000000000016a00000000000000fb3386fd1c",
    x"030b0000000000000155fffffffffffff50003e3ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dd21e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f4ab11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd3a7c1c",
    x"070a0000000000000265fffffffffffff8ef3606841c",
    x"0802000000000000015afffffffffffff6f669ebd81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266e22c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe5911c",
    x"0209000000000000016500000000000000fb3386f81c",
    x"030b0000000000000165fffffffffffff50003e3ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dd21c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f4aad1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd3a761c",
    x"070a000000000000026afffffffffffff8ef3606801c",
    x"080200000000000001a5fffffffffffff6f669ebd51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266e2281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe5931c",
    x"020900000000000002aa00000000000000fb3386f21c",
    x"030b00000000000002aafffffffffffff50003e3ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd21a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f4aa91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd3a701c",
    x"070a0000000000000155fffffffffffff8ef36067d1c",
    x"080200000000000002aafffffffffffff6f669ebd31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e2241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5941c",
    x"0209000000000000031f00000000000000fb3386ed1c",
    x"030b000000000000031ffffffffffffff50003e3f01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd2171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f4aa51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd3a6a1c",
    x"070a000000000000031ffffffffffffff8ef3606791c",
    x"0802000000000000031ffffffffffffff6f669ebd11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e2201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5951c",
    x"020900000000000000ae00000000000000fb3386e71c",
    x"030b00000000000000aefffffffffffff50003e3f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd2151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f4aa21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd3a641c",
    x"070a00000000000000aefffffffffffff8ef3606761c",
    x"080200000000000000aefffffffffffff6f669ebce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e21c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5961c",
    x"020900000000000001a400000000000000fb3386e11c",
    x"030b00000000000001a4fffffffffffff50003e3f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd2131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f4a9e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd3a5d1c",
    x"070a00000000000001a4fffffffffffff8ef3606721c",
    x"080200000000000001a4fffffffffffff6f669ebcc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266e2171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe5971c",
    x"0209000000000000025a00000000000000fb3386dc1c",
    x"030b000000000000025afffffffffffff50003e3f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dd2101c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f4a9a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd3a571c",
    x"070a000000000000025afffffffffffff8ef36066f1c",
    x"0802000000000000025afffffffffffff6f669ebc91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2131c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5981c",
    x"020900000000000002aa00000000000000fb3386d61c",
    x"030b00000000000002aafffffffffffff50003e3f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd20e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a511c",
    x"070a00000000000002aafffffffffffff8ef36066b1c",
    x"080200000000000002aafffffffffffff6f669ebc71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266e20f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe5991c",
    x"0209000000000000029a00000000000000fb3386d11c",
    x"030b000000000000029afffffffffffff50003e3f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dd20c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f4a931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd3a4b1c",
    x"070a000000000000029afffffffffffff8ef3606681c",
    x"0802000000000000029afffffffffffff6f669ebc51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e20b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe59a1c",
    x"020900000000000002aa00000000000000fb3386cb1c",
    x"030b00000000000002aafffffffffffff50003e3f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a8f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a451c",
    x"070a00000000000002aafffffffffffff8ef3606641c",
    x"080200000000000002aafffffffffffff6f669ebc21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe59b1c",
    x"020900000000000002aa00000000000000fb3386c51c",
    x"030b00000000000002aafffffffffffff50003e3f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a8b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a3f1c",
    x"070a00000000000002aafffffffffffff8ef3606601c",
    x"080200000000000002aafffffffffffff6f669ebc01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e2021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe59c1c",
    x"020900000000000002aa00000000000000fb3386c01c",
    x"030b00000000000002aafffffffffffff50003e3f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a391c",
    x"070a00000000000002aafffffffffffff8ef36065d1c",
    x"080200000000000002aafffffffffffff6f669ebbe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1fe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe59d1c",
    x"020900000000000002aa00000000000000fb3386ba1c",
    x"030b00000000000002aafffffffffffff50003e3fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a331c",
    x"070a00000000000002aafffffffffffff8ef3606591c",
    x"080200000000000002aafffffffffffff6f669ebbb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1fa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe59e1c",
    x"020900000000000002aa00000000000000fb3386b51c",
    x"030b00000000000002aafffffffffffff50003e3fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd2001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a2c1c",
    x"070a00000000000002aafffffffffffff8ef3606561c",
    x"080200000000000002aafffffffffffff6f669ebb91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1f61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5a01c",
    x"020900000000000002aa00000000000000fb3386af1c",
    x"030b00000000000002aafffffffffffff50003e3fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1fe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a7c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a261c",
    x"070a00000000000002aafffffffffffff8ef3606521c",
    x"080200000000000002aafffffffffffff6f669ebb61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1f21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5a11c",
    x"020900000000000002aa00000000000000fb3386a91c",
    x"030b00000000000002aafffffffffffff50003e3fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1fb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd3a201c",
    x"070a00000000000002aafffffffffffff8ef36064f1c",
    x"080200000000000002aafffffffffffff6f669ebb41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266e1ed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe5a21c",
    x"0209000000000000016600000000000000fb3386a41c",
    x"030b0000000000000166fffffffffffff50003e3fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dd1f91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f4a751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd3a1a1c",
    x"070a0000000000000166fffffffffffff8ef36064b1c",
    x"08020000000000000166fffffffffffff6f669ebb21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1e91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5a31c",
    x"0209000000000000015500000000000000fb33869e1c",
    x"030b0000000000000155fffffffffffff50003e3ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1f61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a141c",
    x"070a0000000000000155fffffffffffff8ef3606481c",
    x"08020000000000000155fffffffffffff6f669ebaf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1e51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5a41c",
    x"0209000000000000015500000000000000fb3386991c",
    x"030b0000000000000155fffffffffffff50003e4001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1f41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a6d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a0e1c",
    x"070a0000000000000155fffffffffffff8ef3606441c",
    x"08020000000000000155fffffffffffff6f669ebad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1e11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5a51c",
    x"0209000000000000015500000000000000fb3386931c",
    x"030b0000000000000155fffffffffffff50003e4011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1f21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a6a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a081c",
    x"070a0000000000000155fffffffffffff8ef3606411c",
    x"08020000000000000155fffffffffffff6f669ebab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1dd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5a61c",
    x"0209000000000000015500000000000000fb33868e1c",
    x"030b0000000000000155fffffffffffff50003e4021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1ef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd3a021c",
    x"070a0000000000000155fffffffffffff8ef36063d1c",
    x"08020000000000000155fffffffffffff6f669eba81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5a71c",
    x"0209000000000000015500000000000000fb3386881c",
    x"030b0000000000000155fffffffffffff50003e4031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1ed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39fb1c",
    x"070a0000000000000155fffffffffffff8ef3606391c",
    x"08020000000000000155fffffffffffff6f669eba61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266e1d41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe5a81c",
    x"0209000000000000015900000000000000fb3386821c",
    x"030b0000000000000159fffffffffffff50003e4041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dd1eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f4a5e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd39f51c",
    x"070a0000000000000159fffffffffffff8ef3606361c",
    x"08020000000000000159fffffffffffff6f669eba41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e1d01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5a91c",
    x"0209000000000000031f00000000000000fb33867d1c",
    x"030b000000000000031ffffffffffffff50003e4051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd1e81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f4a5b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd39ef1c",
    x"070a000000000000031ffffffffffffff8ef3606321c",
    x"0802000000000000031ffffffffffffff6f669eba11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e1cc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5aa1c",
    x"020900000000000000ae00000000000000fb3386771c",
    x"030b00000000000000aefffffffffffff50003e4061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd1e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f4a571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd39e91c",
    x"070a00000000000000aefffffffffffff8ef36062f1c",
    x"080200000000000000aefffffffffffff6f669eb9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e1c81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5ab1c",
    x"020900000000000001a400000000000000fb3386721c",
    x"030b00000000000001a4fffffffffffff50003e4071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd1e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f4a531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd39e31c",
    x"070a00000000000001a4fffffffffffff8ef36062b1c",
    x"080200000000000001a4fffffffffffff6f669eb9c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266e1c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe5ad1c",
    x"0209000000000000029a00000000000000fb33866c1c",
    x"030b000000000000029afffffffffffff50003e4081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dd1e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f4a4f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd39dd1c",
    x"070a000000000000029afffffffffffff8ef3606281c",
    x"0802000000000000029afffffffffffff6f669eb9a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1bf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5ae1c",
    x"020900000000000002aa00000000000000fb3386661c",
    x"030b00000000000002aafffffffffffff50003e40a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a4c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39d71c",
    x"070a00000000000002aafffffffffffff8ef3606241c",
    x"080200000000000002aafffffffffffff6f669eb981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266e1bb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe5af1c",
    x"0209000000000000029a00000000000000fb3386611c",
    x"030b000000000000029afffffffffffff50003e40b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dd1dd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f4a481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd39d11c",
    x"070a000000000000029afffffffffffff8ef3606211c",
    x"0802000000000000029afffffffffffff6f669eb951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1b71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b01c",
    x"020900000000000002aa00000000000000fb33865b1c",
    x"030b00000000000002aafffffffffffff50003e40c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39ca1c",
    x"070a00000000000002aafffffffffffff8ef36061d1c",
    x"080200000000000002aafffffffffffff6f669eb931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b11c",
    x"020900000000000002aa00000000000000fb3386561c",
    x"030b00000000000002aafffffffffffff50003e40d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1d81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39c41c",
    x"070a00000000000002aafffffffffffff8ef3606191c",
    x"080200000000000002aafffffffffffff6f669eb911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b21c",
    x"020900000000000002aa00000000000000fb3386501c",
    x"030b00000000000002aafffffffffffff50003e40e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1d61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a3d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39be1c",
    x"070a00000000000002aafffffffffffff8ef3606161c",
    x"080200000000000002aafffffffffffff6f669eb8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b31c",
    x"020900000000000002aa00000000000000fb33864b1c",
    x"030b00000000000002aafffffffffffff50003e40f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1d31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39b81c",
    x"070a00000000000002aafffffffffffff8ef3606121c",
    x"080200000000000002aafffffffffffff6f669eb8c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1a61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b41c",
    x"020900000000000002aa00000000000000fb3386451c",
    x"030b00000000000002aafffffffffffff50003e4101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1d11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39b21c",
    x"070a00000000000002aafffffffffffff8ef36060f1c",
    x"080200000000000002aafffffffffffff6f669eb891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b51c",
    x"020900000000000002aa00000000000000fb33863f1c",
    x"030b00000000000002aafffffffffffff50003e4111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1cf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39ac1c",
    x"070a00000000000002aafffffffffffff8ef36060b1c",
    x"080200000000000002aafffffffffffff6f669eb871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e19d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b61c",
    x"020900000000000002aa00000000000000fb33863a1c",
    x"030b00000000000002aafffffffffffff50003e4121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a2e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39a61c",
    x"070a00000000000002aafffffffffffff8ef3606081c",
    x"080200000000000002aafffffffffffff6f669eb851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b71c",
    x"020900000000000002aa00000000000000fb3386341c",
    x"030b00000000000002aafffffffffffff50003e4131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1ca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a2a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39a01c",
    x"070a00000000000002aafffffffffffff8ef3606041c",
    x"080200000000000002aafffffffffffff6f669eb821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5b91c",
    x"020900000000000002aa00000000000000fb33862f1c",
    x"030b00000000000002aafffffffffffff50003e4141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1c81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a261c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39991c",
    x"070a00000000000002aafffffffffffff8ef3606011c",
    x"080200000000000002aafffffffffffff6f669eb801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5ba1c",
    x"020900000000000002aa00000000000000fb3386291c",
    x"030b00000000000002aafffffffffffff50003e4151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39931c",
    x"070a00000000000002aafffffffffffff8ef3605fd1c",
    x"080200000000000002aafffffffffffff6f669eb7e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e18d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5bb1c",
    x"020900000000000002aa00000000000000fb3386231c",
    x"030b00000000000002aafffffffffffff50003e4161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1c31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a1f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd398d1c",
    x"070a00000000000002aafffffffffffff8ef3605fa1c",
    x"080200000000000002aafffffffffffff6f669eb7b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e1881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5bc1c",
    x"020900000000000002aa00000000000000fb33861e1c",
    x"030b00000000000002aafffffffffffff50003e4171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1c11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f4a1b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd39871c",
    x"070a00000000000002aafffffffffffff8ef3605f61c",
    x"080200000000000002aafffffffffffff6f669eb791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266e1841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbe5bd1c",
    x"020900000000000001aa00000000000000fb3386181c",
    x"030b00000000000001aafffffffffffff50003e4181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dd1be1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f4a171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd39811c",
    x"070a00000000000001aafffffffffffff8ef3605f21c",
    x"080200000000000001aafffffffffffff6f669eb771c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5be1c",
    x"0209000000000000015500000000000000fb3386131c",
    x"030b0000000000000155fffffffffffff50003e4191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1bc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd397b1c",
    x"070a0000000000000155fffffffffffff8ef3605ef1c",
    x"08020000000000000155fffffffffffff6f669eb741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e17c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5bf1c",
    x"0209000000000000031f00000000000000fb33860d1c",
    x"030b000000000000031ffffffffffffff50003e41a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd1b91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f4a101c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd39751c",
    x"070a000000000000031ffffffffffffff8ef3605eb1c",
    x"0802000000000000031ffffffffffffff6f669eb721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e1781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5c01c",
    x"020900000000000000ae00000000000000fb3386071c",
    x"030b00000000000000aefffffffffffff50003e41b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd1b71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f4a0c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd396f1c",
    x"070a00000000000000aefffffffffffff8ef3605e81c",
    x"080200000000000000aefffffffffffff6f669eb6f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e1731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5c11c",
    x"020900000000000001a400000000000000fb3386021c",
    x"030b00000000000001a4fffffffffffff50003e41c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd1b51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f4a081c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd39681c",
    x"070a00000000000001a4fffffffffffff8ef3605e41c",
    x"080200000000000001a4fffffffffffff6f669eb6d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266e16f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe5c21c",
    x"0209000000000000019a00000000000000fb3385fc1c",
    x"030b000000000000019afffffffffffff50003e41e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dd1b21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f4a051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd39621c",
    x"070a000000000000019afffffffffffff8ef3605e11c",
    x"0802000000000000019afffffffffffff6f669eb6b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e16b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5c31c",
    x"0209000000000000015500000000000000fb3385f71c",
    x"030b0000000000000155fffffffffffff50003e41f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1b01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f4a011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd395c1c",
    x"070a0000000000000155fffffffffffff8ef3605dd1c",
    x"08020000000000000155fffffffffffff6f669eb681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5c41c",
    x"0209000000000000015500000000000000fb3385f11c",
    x"030b0000000000000155fffffffffffff50003e4201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49fd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39561c",
    x"070a0000000000000155fffffffffffff8ef3605da1c",
    x"08020000000000000155fffffffffffff6f669eb661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5c61c",
    x"0209000000000000015500000000000000fb3385ec1c",
    x"030b0000000000000155fffffffffffff50003e4211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1ab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49fa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39501c",
    x"070a0000000000000155fffffffffffff8ef3605d61c",
    x"08020000000000000155fffffffffffff6f669eb641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e15e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5c71c",
    x"0209000000000000015500000000000000fb3385e61c",
    x"030b0000000000000155fffffffffffff50003e4221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49f61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd394a1c",
    x"070a0000000000000155fffffffffffff8ef3605d21c",
    x"08020000000000000155fffffffffffff6f669eb611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e15a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5c81c",
    x"0209000000000000015500000000000000fb3385e01c",
    x"030b0000000000000155fffffffffffff50003e4231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1a71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49f21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39441c",
    x"070a0000000000000155fffffffffffff8ef3605cf1c",
    x"08020000000000000155fffffffffffff6f669eb5f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5c91c",
    x"0209000000000000015500000000000000fb3385db1c",
    x"030b0000000000000155fffffffffffff50003e4241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49ee1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd393d1c",
    x"070a0000000000000155fffffffffffff8ef3605cb1c",
    x"08020000000000000155fffffffffffff6f669eb5c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5ca1c",
    x"0209000000000000015500000000000000fb3385d51c",
    x"030b0000000000000155fffffffffffff50003e4251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39371c",
    x"070a0000000000000155fffffffffffff8ef3605c81c",
    x"08020000000000000155fffffffffffff6f669eb5a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e14e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5cb1c",
    x"0209000000000000015500000000000000fb3385d01c",
    x"030b0000000000000155fffffffffffff50003e4261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1a01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49e71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39311c",
    x"070a0000000000000155fffffffffffff8ef3605c41c",
    x"08020000000000000155fffffffffffff6f669eb581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1491c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5cc1c",
    x"0209000000000000015500000000000000fb3385ca1c",
    x"030b0000000000000155fffffffffffff50003e4271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd19d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49e31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd392b1c",
    x"070a0000000000000155fffffffffffff8ef3605c11c",
    x"08020000000000000155fffffffffffff6f669eb551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1451c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5cd1c",
    x"0209000000000000015500000000000000fb3385c41c",
    x"030b0000000000000155fffffffffffff50003e4281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd19b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49df1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39251c",
    x"070a0000000000000155fffffffffffff8ef3605bd1c",
    x"08020000000000000155fffffffffffff6f669eb531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1411c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5ce1c",
    x"0209000000000000015500000000000000fb3385bf1c",
    x"030b0000000000000155fffffffffffff50003e4291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1991c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49dc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd391f1c",
    x"070a0000000000000155fffffffffffff8ef3605ba1c",
    x"08020000000000000155fffffffffffff6f669eb511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e13d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5cf1c",
    x"0209000000000000015500000000000000fb3385b91c",
    x"030b0000000000000155fffffffffffff50003e42a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49d81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39191c",
    x"070a0000000000000155fffffffffffff8ef3605b61c",
    x"08020000000000000155fffffffffffff6f669eb4e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5d01c",
    x"0209000000000000015500000000000000fb3385b41c",
    x"030b0000000000000155fffffffffffff50003e42b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1941c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49d41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39131c",
    x"070a0000000000000155fffffffffffff8ef3605b21c",
    x"08020000000000000155fffffffffffff6f669eb4c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5d21c",
    x"0209000000000000015500000000000000fb3385ae1c",
    x"030b0000000000000155fffffffffffff50003e42c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd390c1c",
    x"070a0000000000000155fffffffffffff8ef3605af1c",
    x"08020000000000000155fffffffffffff6f669eb491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5d31c",
    x"0209000000000000015500000000000000fb3385a91c",
    x"030b0000000000000155fffffffffffff50003e42d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd18f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49cd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39061c",
    x"070a0000000000000155fffffffffffff8ef3605ab1c",
    x"08020000000000000155fffffffffffff6f669eb471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e12c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5d41c",
    x"0209000000000000015500000000000000fb3385a31c",
    x"030b0000000000000155fffffffffffff50003e42e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd18d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd39001c",
    x"070a0000000000000155fffffffffffff8ef3605a81c",
    x"08020000000000000155fffffffffffff6f669eb451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e1281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5d51c",
    x"0209000000000000031f00000000000000fb33859d1c",
    x"030b000000000000031ffffffffffffff50003e42f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd18a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f49c51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd38fa1c",
    x"070a000000000000031ffffffffffffff8ef3605a41c",
    x"0802000000000000031ffffffffffffff6f669eb421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e1231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5d61c",
    x"020900000000000000ae00000000000000fb3385981c",
    x"030b00000000000000aefffffffffffff50003e4301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd1881c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f49c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd38f41c",
    x"070a00000000000000aefffffffffffff8ef3605a11c",
    x"080200000000000000aefffffffffffff6f669eb401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e11f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5d71c",
    x"020900000000000001a400000000000000fb3385921c",
    x"030b00000000000001a4fffffffffffff50003e4311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd1861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f49be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd38ee1c",
    x"070a00000000000001a4fffffffffffff8ef36059d1c",
    x"080200000000000001a4fffffffffffff6f669eb3e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266e11b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe5d81c",
    x"0209000000000000015600000000000000fb33858d1c",
    x"030b0000000000000156fffffffffffff50003e4321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dd1831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f49ba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd38e81c",
    x"070a0000000000000156fffffffffffff8ef36059a1c",
    x"08020000000000000156fffffffffffff6f669eb3b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266e1171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe5d91c",
    x"0209000000000000029500000000000000fb3385871c",
    x"030b0000000000000295fffffffffffff50003e4341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd1811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f49b61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd38e21c",
    x"070a0000000000000295fffffffffffff8ef3605961c",
    x"08020000000000000295fffffffffffff6f669eb391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1131c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5da1c",
    x"0209000000000000015500000000000000fb3385811c",
    x"030b0000000000000155fffffffffffff50003e4351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd17f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38db1c",
    x"070a0000000000000155fffffffffffff8ef3605921c",
    x"08020000000000000155fffffffffffff6f669eb371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e10e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5db1c",
    x"0209000000000000015500000000000000fb33857c1c",
    x"030b0000000000000155fffffffffffff50003e4361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd17c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49af1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38d51c",
    x"070a0000000000000155fffffffffffff8ef36058f1c",
    x"08020000000000000155fffffffffffff6f669eb341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e10a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5dc1c",
    x"0209000000000000015500000000000000fb3385761c",
    x"030b0000000000000155fffffffffffff50003e4371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd17a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49ab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38cf1c",
    x"070a0000000000000155fffffffffffff8ef36058b1c",
    x"08020000000000000155fffffffffffff6f669eb321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5dd1c",
    x"0209000000000000015500000000000000fb3385711c",
    x"030b0000000000000155fffffffffffff50003e4381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49a71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38c91c",
    x"070a0000000000000155fffffffffffff8ef3605881c",
    x"08020000000000000155fffffffffffff6f669eb2f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e1021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5df1c",
    x"0209000000000000015500000000000000fb33856b1c",
    x"030b0000000000000155fffffffffffff50003e4391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49a41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38c31c",
    x"070a0000000000000155fffffffffffff8ef3605841c",
    x"08020000000000000155fffffffffffff6f669eb2d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0fe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e01c",
    x"0209000000000000015500000000000000fb3385651c",
    x"030b0000000000000155fffffffffffff50003e43a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49a01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38bd1c",
    x"070a0000000000000155fffffffffffff8ef3605811c",
    x"08020000000000000155fffffffffffff6f669eb2b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e11c",
    x"0209000000000000015500000000000000fb3385601c",
    x"030b0000000000000155fffffffffffff50003e43b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f499c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38b71c",
    x"070a0000000000000155fffffffffffff8ef36057d1c",
    x"08020000000000000155fffffffffffff6f669eb281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e21c",
    x"0209000000000000015500000000000000fb33855a1c",
    x"030b0000000000000155fffffffffffff50003e43c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd16e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49991c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38b11c",
    x"070a0000000000000155fffffffffffff8ef36057a1c",
    x"08020000000000000155fffffffffffff6f669eb261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0f11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e31c",
    x"0209000000000000015500000000000000fb3385551c",
    x"030b0000000000000155fffffffffffff50003e43d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd16c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49951c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38aa1c",
    x"070a0000000000000155fffffffffffff8ef3605761c",
    x"08020000000000000155fffffffffffff6f669eb241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0ed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e41c",
    x"0209000000000000015500000000000000fb33854f1c",
    x"030b0000000000000155fffffffffffff50003e43e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd16a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38a41c",
    x"070a0000000000000155fffffffffffff8ef3605721c",
    x"08020000000000000155fffffffffffff6f669eb211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0e91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e51c",
    x"0209000000000000015500000000000000fb33854a1c",
    x"030b0000000000000155fffffffffffff50003e43f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f498d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd389e1c",
    x"070a0000000000000155fffffffffffff8ef36056f1c",
    x"08020000000000000155fffffffffffff6f669eb1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e61c",
    x"0209000000000000015500000000000000fb3385441c",
    x"030b0000000000000155fffffffffffff50003e4401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f498a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38981c",
    x"070a0000000000000155fffffffffffff8ef36056b1c",
    x"08020000000000000155fffffffffffff6f669eb1c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe5e71c",
    x"0209000000000000015500000000000000fb33853e1c",
    x"030b0000000000000155fffffffffffff50003e4411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1621c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd38921c",
    x"070a0000000000000155fffffffffffff8ef3605681c",
    x"08020000000000000155fffffffffffff6f669eb1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266e0dc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe5e81c",
    x"0209000000000000019500000000000000fb3385391c",
    x"030b0000000000000195fffffffffffff50003e4421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dd1601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f49821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000195ffffffffffffff04cd388c1c",
    x"070a0000000000000195fffffffffffff8ef3605641c",
    x"08020000000000000195fffffffffffff6f669eb181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5e91c",
    x"020900000000000002aa00000000000000fb3385331c",
    x"030b00000000000002aafffffffffffff50003e4431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd15e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f497e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38861c",
    x"070a00000000000002aafffffffffffff8ef3605611c",
    x"080200000000000002aafffffffffffff6f669eb151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e0d41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe5eb1c",
    x"0209000000000000031f00000000000000fb33852e1c",
    x"030b000000000000031ffffffffffffff50003e4441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd15b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f497b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd387f1c",
    x"070a000000000000031ffffffffffffff8ef36055d1c",
    x"0802000000000000031ffffffffffffff6f669eb131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e0cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe5ec1c",
    x"020900000000000000ae00000000000000fb3385281c",
    x"030b00000000000000aefffffffffffff50003e4451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd1591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f49771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd38791c",
    x"070a00000000000000aefffffffffffff8ef36055a1c",
    x"080200000000000000aefffffffffffff6f669eb111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e0cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe5ed1c",
    x"020900000000000001a400000000000000fb3385221c",
    x"030b00000000000001a4fffffffffffff50003e4461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd1571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f49731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd38731c",
    x"070a00000000000001a4fffffffffffff8ef3605561c",
    x"080200000000000001a4fffffffffffff6f669eb0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266e0c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe5ee1c",
    x"0209000000000000025600000000000000fb33851d1c",
    x"030b0000000000000256fffffffffffff50003e4471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dd1541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f496f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd386d1c",
    x"070a0000000000000256fffffffffffff8ef3605521c",
    x"08020000000000000256fffffffffffff6f669eb0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5ef1c",
    x"020900000000000002aa00000000000000fb3385171c",
    x"030b00000000000002aafffffffffffff50003e4481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f496c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38671c",
    x"070a00000000000002aafffffffffffff8ef36054f1c",
    x"080200000000000002aafffffffffffff6f669eb091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0bf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f01c",
    x"020900000000000002aa00000000000000fb3385121c",
    x"030b00000000000002aafffffffffffff50003e44a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38611c",
    x"070a00000000000002aafffffffffffff8ef36054b1c",
    x"080200000000000002aafffffffffffff6f669eb071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f11c",
    x"020900000000000002aa00000000000000fb33850c1c",
    x"030b00000000000002aafffffffffffff50003e44b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd14d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd385b1c",
    x"070a00000000000002aafffffffffffff8ef3605481c",
    x"080200000000000002aafffffffffffff6f669eb051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f21c",
    x"020900000000000002aa00000000000000fb3385061c",
    x"030b00000000000002aafffffffffffff50003e44c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd14b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38551c",
    x"070a00000000000002aafffffffffffff8ef3605441c",
    x"080200000000000002aafffffffffffff6f669eb021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f31c",
    x"020900000000000002aa00000000000000fb3385011c",
    x"030b00000000000002aafffffffffffff50003e44d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f495d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd384e1c",
    x"070a00000000000002aafffffffffffff8ef3605411c",
    x"080200000000000002aafffffffffffff6f669eb001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f41c",
    x"020900000000000002aa00000000000000fb3384fb1c",
    x"030b00000000000002aafffffffffffff50003e44e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38481c",
    x"070a00000000000002aafffffffffffff8ef36053d1c",
    x"080200000000000002aafffffffffffff6f669eafe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f51c",
    x"020900000000000002aa00000000000000fb3384f61c",
    x"030b00000000000002aafffffffffffff50003e44f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38421c",
    x"070a00000000000002aafffffffffffff8ef36053a1c",
    x"080200000000000002aafffffffffffff6f669eafb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f61c",
    x"020900000000000002aa00000000000000fb3384f01c",
    x"030b00000000000002aafffffffffffff50003e4501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd383c1c",
    x"070a00000000000002aafffffffffffff8ef3605361c",
    x"080200000000000002aafffffffffffff6f669eaf91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f81c",
    x"020900000000000002aa00000000000000fb3384eb1c",
    x"030b00000000000002aafffffffffffff50003e4511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd13f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f494e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38361c",
    x"070a00000000000002aafffffffffffff8ef3605321c",
    x"080200000000000002aafffffffffffff6f669eaf71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e09d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5f91c",
    x"020900000000000002aa00000000000000fb3384e51c",
    x"030b00000000000002aafffffffffffff50003e4521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd13d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f494a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38301c",
    x"070a00000000000002aafffffffffffff8ef36052f1c",
    x"080200000000000002aafffffffffffff6f669eaf41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5fa1c",
    x"020900000000000002aa00000000000000fb3384df1c",
    x"030b00000000000002aafffffffffffff50003e4531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd13a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49461c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd382a1c",
    x"070a00000000000002aafffffffffffff8ef36052b1c",
    x"080200000000000002aafffffffffffff6f669eaf21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5fb1c",
    x"020900000000000002aa00000000000000fb3384da1c",
    x"030b00000000000002aafffffffffffff50003e4541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49431c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38241c",
    x"070a00000000000002aafffffffffffff8ef3605281c",
    x"080200000000000002aafffffffffffff6f669eaef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5fc1c",
    x"020900000000000002aa00000000000000fb3384d41c",
    x"030b00000000000002aafffffffffffff50003e4551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f493f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd381d1c",
    x"070a00000000000002aafffffffffffff8ef3605241c",
    x"080200000000000002aafffffffffffff6f669eaed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e08c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5fd1c",
    x"020900000000000002aa00000000000000fb3384cf1c",
    x"030b00000000000002aafffffffffffff50003e4561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f493b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd38171c",
    x"070a00000000000002aafffffffffffff8ef3605211c",
    x"080200000000000002aafffffffffffff6f669eaeb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266e0881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe5fe1c",
    x"0209000000000000029a00000000000000fb3384c91c",
    x"030b000000000000029afffffffffffff50003e4571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dd1311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f49381c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd38111c",
    x"070a000000000000029afffffffffffff8ef36051d1c",
    x"0802000000000000029afffffffffffff6f669eae81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e0841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe5ff1c",
    x"020900000000000002aa00000000000000fb3384c31c",
    x"030b00000000000002aafffffffffffff50003e4581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd12f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd380b1c",
    x"070a00000000000002aafffffffffffff8ef36051a1c",
    x"080200000000000002aafffffffffffff6f669eae61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e0801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6001c",
    x"0209000000000000031f00000000000000fb3384be1c",
    x"030b000000000000031ffffffffffffff50003e4591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd12c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f49301c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd38051c",
    x"070a000000000000031ffffffffffffff8ef3605161c",
    x"0802000000000000031ffffffffffffff6f669eae41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e07b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6011c",
    x"020900000000000000ae00000000000000fb3384b81c",
    x"030b00000000000000aefffffffffffff50003e45a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd12a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f492c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd37ff1c",
    x"070a00000000000000aefffffffffffff8ef3605121c",
    x"080200000000000000aefffffffffffff6f669eae11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e0771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6021c",
    x"020900000000000001a400000000000000fb3384b31c",
    x"030b00000000000001a4fffffffffffff50003e45b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd1281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f49291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd37f91c",
    x"070a00000000000001a4fffffffffffff8ef36050f1c",
    x"080200000000000001a4fffffffffffff6f669eadf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266e0731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe6041c",
    x"0209000000000000029600000000000000fb3384ad1c",
    x"030b0000000000000296fffffffffffff50003e45c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dd1251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f49251c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd37f31c",
    x"070a0000000000000296fffffffffffff8ef36050b1c",
    x"08020000000000000296fffffffffffff6f669eadc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266e06f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6051c",
    x"020900000000000002aa00000000000000fb3384a71c",
    x"030b00000000000002aafffffffffffff50003e45d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd1231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f49211c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd37ec1c",
    x"070a00000000000002aafffffffffffff8ef3605081c",
    x"080200000000000002aafffffffffffff6f669eada1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266e06a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe6061c",
    x"0209000000000000016500000000000000fb3384a21c",
    x"030b0000000000000165fffffffffffff50003e45e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dd1211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f491d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd37e61c",
    x"070a0000000000000165fffffffffffff8ef3605041c",
    x"08020000000000000165fffffffffffff6f669ead81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6071c",
    x"0209000000000000015500000000000000fb33849c1c",
    x"030b0000000000000155fffffffffffff50003e45f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd11e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f491a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37e01c",
    x"070a0000000000000155fffffffffffff8ef3605011c",
    x"08020000000000000155fffffffffffff6f669ead51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6081c",
    x"0209000000000000015500000000000000fb3384971c",
    x"030b0000000000000155fffffffffffff50003e4601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd11c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49161c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37da1c",
    x"070a0000000000000155fffffffffffff8ef3604fd1c",
    x"08020000000000000155fffffffffffff6f669ead31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e05e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6091c",
    x"0209000000000000015500000000000000fb3384911c",
    x"030b0000000000000155fffffffffffff50003e4621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37d41c",
    x"070a0000000000000155fffffffffffff8ef3604fa1c",
    x"08020000000000000155fffffffffffff6f669ead11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e05a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe60a1c",
    x"0209000000000000015500000000000000fb33848c1c",
    x"030b0000000000000155fffffffffffff50003e4631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f490f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37ce1c",
    x"070a0000000000000155fffffffffffff8ef3604f61c",
    x"08020000000000000155fffffffffffff6f669eace1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe60b1c",
    x"0209000000000000015500000000000000fb3384861c",
    x"030b0000000000000155fffffffffffff50003e4641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f490b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37c81c",
    x"070a0000000000000155fffffffffffff8ef3604f21c",
    x"08020000000000000155fffffffffffff6f669eacc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe60c1c",
    x"0209000000000000015500000000000000fb3384801c",
    x"030b0000000000000155fffffffffffff50003e4651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37c11c",
    x"070a0000000000000155fffffffffffff8ef3604ef1c",
    x"08020000000000000155fffffffffffff6f669eac91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e04d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe60d1c",
    x"0209000000000000015500000000000000fb33847b1c",
    x"030b0000000000000155fffffffffffff50003e4661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1101c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37bb1c",
    x"070a0000000000000155fffffffffffff8ef3604eb1c",
    x"08020000000000000155fffffffffffff6f669eac71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0491c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe60e1c",
    x"0209000000000000015500000000000000fb3384751c",
    x"030b0000000000000155fffffffffffff50003e4671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd10e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f49001c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37b51c",
    x"070a0000000000000155fffffffffffff8ef3604e81c",
    x"08020000000000000155fffffffffffff6f669eac51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0451c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6101c",
    x"0209000000000000015500000000000000fb3384701c",
    x"030b0000000000000155fffffffffffff50003e4681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd10b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48fc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37af1c",
    x"070a0000000000000155fffffffffffff8ef3604e41c",
    x"08020000000000000155fffffffffffff6f669eac21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6111c",
    x"0209000000000000015500000000000000fb33846a1c",
    x"030b0000000000000155fffffffffffff50003e4691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37a91c",
    x"070a0000000000000155fffffffffffff8ef3604e11c",
    x"08020000000000000155fffffffffffff6f669eac01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e03c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6121c",
    x"0209000000000000015500000000000000fb3384641c",
    x"030b0000000000000155fffffffffffff50003e46a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37a31c",
    x"070a0000000000000155fffffffffffff8ef3604dd1c",
    x"08020000000000000155fffffffffffff6f669eabe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6131c",
    x"0209000000000000015500000000000000fb33845f1c",
    x"030b0000000000000155fffffffffffff50003e46b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48f11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd379d1c",
    x"070a0000000000000155fffffffffffff8ef3604d91c",
    x"08020000000000000155fffffffffffff6f669eabb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266e0341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe6141c",
    x"0209000000000000025500000000000000fb3384591c",
    x"030b0000000000000255fffffffffffff50003e46c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dd1021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f48ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd37971c",
    x"070a0000000000000255fffffffffffff8ef3604d61c",
    x"08020000000000000255fffffffffffff6f669eab91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6151c",
    x"0209000000000000015500000000000000fb3384541c",
    x"030b0000000000000155fffffffffffff50003e46d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd1001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37901c",
    x"070a0000000000000155fffffffffffff8ef3604d21c",
    x"08020000000000000155fffffffffffff6f669eab61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266e02b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6161c",
    x"0209000000000000031f00000000000000fb33844e1c",
    x"030b000000000000031ffffffffffffff50003e46e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd0fd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f48e61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd378a1c",
    x"070a000000000000031ffffffffffffff8ef3604cf1c",
    x"0802000000000000031ffffffffffffff6f669eab41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266e0271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6171c",
    x"020900000000000000ae00000000000000fb3384491c",
    x"030b00000000000000aefffffffffffff50003e46f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd0fb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f48e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd37841c",
    x"070a00000000000000aefffffffffffff8ef3604cb1c",
    x"080200000000000000aefffffffffffff6f669eab21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266e0231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6181c",
    x"020900000000000001a400000000000000fb3384431c",
    x"030b00000000000001a4fffffffffffff50003e4701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd0f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f48de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd377e1c",
    x"070a00000000000001a4fffffffffffff8ef3604c81c",
    x"080200000000000001a4fffffffffffff6f669eaaf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266e01f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe6191c",
    x"0209000000000000019600000000000000fb33843d1c",
    x"030b0000000000000196fffffffffffff50003e4711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dd0f61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f48da1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000196ffffffffffffff04cd37781c",
    x"070a0000000000000196fffffffffffff8ef3604c41c",
    x"08020000000000000196fffffffffffff6f669eaad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e01b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe61a1c",
    x"0209000000000000015500000000000000fb3384381c",
    x"030b0000000000000155fffffffffffff50003e4721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0f41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48d71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37721c",
    x"070a0000000000000155fffffffffffff8ef3604c11c",
    x"08020000000000000155fffffffffffff6f669eaab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe61b1c",
    x"0209000000000000015500000000000000fb3384321c",
    x"030b0000000000000155fffffffffffff50003e4731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0f11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48d31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd376c1c",
    x"070a0000000000000155fffffffffffff8ef3604bd1c",
    x"08020000000000000155fffffffffffff6f669eaa81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe61d1c",
    x"0209000000000000015500000000000000fb33842d1c",
    x"030b0000000000000155fffffffffffff50003e4741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0ef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48cf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37661c",
    x"070a0000000000000155fffffffffffff8ef3604b91c",
    x"08020000000000000155fffffffffffff6f669eaa61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e00e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe61e1c",
    x"0209000000000000015500000000000000fb3384271c",
    x"030b0000000000000155fffffffffffff50003e4751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0ed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48cb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd375f1c",
    x"070a0000000000000155fffffffffffff8ef3604b61c",
    x"08020000000000000155fffffffffffff6f669eaa41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e00a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe61f1c",
    x"0209000000000000015500000000000000fb3384211c",
    x"030b0000000000000155fffffffffffff50003e4761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0ea1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48c81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37591c",
    x"070a0000000000000155fffffffffffff8ef3604b21c",
    x"08020000000000000155fffffffffffff6f669eaa11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6201c",
    x"0209000000000000015500000000000000fb33841c1c",
    x"030b0000000000000155fffffffffffff50003e4771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0e81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48c41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37531c",
    x"070a0000000000000155fffffffffffff8ef3604af1c",
    x"08020000000000000155fffffffffffff6f669ea9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266e0011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6211c",
    x"0209000000000000015500000000000000fb3384161c",
    x"030b0000000000000155fffffffffffff50003e4781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48c01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd374d1c",
    x"070a0000000000000155fffffffffffff8ef3604ab1c",
    x"08020000000000000155fffffffffffff6f669ea9c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dffd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6221c",
    x"0209000000000000015500000000000000fb3384111c",
    x"030b0000000000000155fffffffffffff50003e4791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0e31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48bd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37471c",
    x"070a0000000000000155fffffffffffff8ef3604a81c",
    x"08020000000000000155fffffffffffff6f669ea9a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dff91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6231c",
    x"0209000000000000015500000000000000fb33840b1c",
    x"030b0000000000000155fffffffffffff50003e47b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48b91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37411c",
    x"070a0000000000000155fffffffffffff8ef3604a41c",
    x"08020000000000000155fffffffffffff6f669ea981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dff51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6241c",
    x"0209000000000000015500000000000000fb3384051c",
    x"030b0000000000000155fffffffffffff50003e47c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48b51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd373b1c",
    x"070a0000000000000155fffffffffffff8ef3604a11c",
    x"08020000000000000155fffffffffffff6f669ea951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dff11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6251c",
    x"0209000000000000015500000000000000fb3384001c",
    x"030b0000000000000155fffffffffffff50003e47d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0dc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48b11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37341c",
    x"070a0000000000000155fffffffffffff8ef36049d1c",
    x"08020000000000000155fffffffffffff6f669ea931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6261c",
    x"0209000000000000015500000000000000fb3383fa1c",
    x"030b0000000000000155fffffffffffff50003e47e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48ae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd372e1c",
    x"070a0000000000000155fffffffffffff8ef3604991c",
    x"08020000000000000155fffffffffffff6f669ea911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfe81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6271c",
    x"0209000000000000015500000000000000fb3383f51c",
    x"030b0000000000000155fffffffffffff50003e47f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0d71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48aa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37281c",
    x"070a0000000000000155fffffffffffff8ef3604961c",
    x"08020000000000000155fffffffffffff6f669ea8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfe41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6291c",
    x"0209000000000000015500000000000000fb3383ef1c",
    x"030b0000000000000155fffffffffffff50003e4801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0d51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48a61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd37221c",
    x"070a0000000000000155fffffffffffff8ef3604921c",
    x"08020000000000000155fffffffffffff6f669ea8c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266dfe01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbe62a1c",
    x"020900000000000002a500000000000000fb3383e91c",
    x"030b00000000000002a5fffffffffffff50003e4811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dd0d31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f48a21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd371c1c",
    x"070a00000000000002a5fffffffffffff8ef36048f1c",
    x"080200000000000002a5fffffffffffff6f669ea891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dfdc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe62b1c",
    x"020900000000000002aa00000000000000fb3383e41c",
    x"030b00000000000002aafffffffffffff50003e4821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0d01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f489f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd37161c",
    x"070a00000000000002aafffffffffffff8ef36048b1c",
    x"080200000000000002aafffffffffffff6f669ea871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dfd71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe62c1c",
    x"0209000000000000031f00000000000000fb3383de1c",
    x"030b000000000000031ffffffffffffff50003e4831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd0ce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f489b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd37101c",
    x"070a000000000000031ffffffffffffff8ef3604881c",
    x"0802000000000000031ffffffffffffff6f669ea851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dfd31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe62d1c",
    x"020900000000000000ae00000000000000fb3383d91c",
    x"030b00000000000000aefffffffffffff50003e4841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd0cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f48971c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd370a1c",
    x"070a00000000000000aefffffffffffff8ef3604841c",
    x"080200000000000000aefffffffffffff6f669ea821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dfcf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe62e1c",
    x"020900000000000001a400000000000000fb3383d31c",
    x"030b00000000000001a4fffffffffffff50003e4851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd0c91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f48941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd37031c",
    x"070a00000000000001a4fffffffffffff8ef3604801c",
    x"080200000000000001a4fffffffffffff6f669ea801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266dfcb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbe62f1c",
    x"020900000000000002a600000000000000fb3383ce1c",
    x"030b00000000000002a6fffffffffffff50003e4861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dd0c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f48901c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd36fd1c",
    x"070a00000000000002a6fffffffffffff8ef36047d1c",
    x"080200000000000002a6fffffffffffff6f669ea7e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dfc71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6301c",
    x"020900000000000002aa00000000000000fb3383c81c",
    x"030b00000000000002aafffffffffffff50003e4871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f488c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd36f71c",
    x"070a00000000000002aafffffffffffff8ef3604791c",
    x"080200000000000002aafffffffffffff6f669ea7b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266dfc21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe6311c",
    x"0209000000000000016900000000000000fb3383c21c",
    x"030b0000000000000169fffffffffffff50003e4881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dd0c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001690000000000000b072f48881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd36f11c",
    x"070a0000000000000169fffffffffffff8ef3604761c",
    x"08020000000000000169fffffffffffff6f669ea791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfbe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6321c",
    x"0209000000000000015500000000000000fb3383bd1c",
    x"030b0000000000000155fffffffffffff50003e4891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0c01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48851c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36eb1c",
    x"070a0000000000000155fffffffffffff8ef3604721c",
    x"08020000000000000155fffffffffffff6f669ea761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6331c",
    x"0209000000000000015500000000000000fb3383b71c",
    x"030b0000000000000155fffffffffffff50003e48a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48811c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36e51c",
    x"070a0000000000000155fffffffffffff8ef36046f1c",
    x"08020000000000000155fffffffffffff6f669ea741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfb61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6351c",
    x"0209000000000000015500000000000000fb3383b21c",
    x"030b0000000000000155fffffffffffff50003e48b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f487d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36df1c",
    x"070a0000000000000155fffffffffffff8ef36046b1c",
    x"08020000000000000155fffffffffffff6f669ea721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfb21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6361c",
    x"0209000000000000015500000000000000fb3383ac1c",
    x"030b0000000000000155fffffffffffff50003e48c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0b91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36d81c",
    x"070a0000000000000155fffffffffffff8ef3604681c",
    x"08020000000000000155fffffffffffff6f669ea6f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6371c",
    x"0209000000000000015500000000000000fb3383a61c",
    x"030b0000000000000155fffffffffffff50003e48d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36d21c",
    x"070a0000000000000155fffffffffffff8ef3604641c",
    x"08020000000000000155fffffffffffff6f669ea6d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfa91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6381c",
    x"0209000000000000015500000000000000fb3383a11c",
    x"030b0000000000000155fffffffffffff50003e48e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0b41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36cc1c",
    x"070a0000000000000155fffffffffffff8ef3604601c",
    x"08020000000000000155fffffffffffff6f669ea6b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfa51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6391c",
    x"0209000000000000015500000000000000fb33839b1c",
    x"030b0000000000000155fffffffffffff50003e48f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0b21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f486e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36c61c",
    x"070a0000000000000155fffffffffffff8ef36045d1c",
    x"08020000000000000155fffffffffffff6f669ea681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dfa11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe63a1c",
    x"0209000000000000015500000000000000fb3383961c",
    x"030b0000000000000155fffffffffffff50003e4901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0af1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f486b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36c01c",
    x"070a0000000000000155fffffffffffff8ef3604591c",
    x"08020000000000000155fffffffffffff6f669ea661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df9d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe63b1c",
    x"0209000000000000015500000000000000fb3383901c",
    x"030b0000000000000155fffffffffffff50003e4911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0ad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36ba1c",
    x"070a0000000000000155fffffffffffff8ef3604561c",
    x"08020000000000000155fffffffffffff6f669ea631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe63c1c",
    x"0209000000000000015500000000000000fb33838a1c",
    x"030b0000000000000155fffffffffffff50003e4921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0ab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48631c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36b41c",
    x"070a0000000000000155fffffffffffff8ef3604521c",
    x"08020000000000000155fffffffffffff6f669ea611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe63d1c",
    x"0209000000000000015500000000000000fb3383851c",
    x"030b0000000000000155fffffffffffff50003e4931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0a81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f485f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36ae1c",
    x"070a0000000000000155fffffffffffff8ef36044f1c",
    x"08020000000000000155fffffffffffff6f669ea5f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe63e1c",
    x"0209000000000000015500000000000000fb33837f1c",
    x"030b0000000000000155fffffffffffff50003e4951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0a61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f485c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36a71c",
    x"070a0000000000000155fffffffffffff8ef36044b1c",
    x"08020000000000000155fffffffffffff6f669ea5c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266df8c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe63f1c",
    x"0209000000000000019500000000000000fb33837a1c",
    x"030b0000000000000195fffffffffffff50003e4961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dd0a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f48581c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000195ffffffffffffff04cd36a11c",
    x"070a0000000000000195fffffffffffff8ef3604471c",
    x"08020000000000000195fffffffffffff6f669ea5a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266df881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6411c",
    x"020900000000000002aa00000000000000fb3383741c",
    x"030b00000000000002aafffffffffffff50003e4971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0a11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f48541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd369b1c",
    x"070a00000000000002aafffffffffffff8ef3604441c",
    x"080200000000000002aafffffffffffff6f669ea581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266df831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6421c",
    x"0209000000000000031f00000000000000fb33836f1c",
    x"030b000000000000031ffffffffffffff50003e4981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd09f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f48511c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd36951c",
    x"070a000000000000031ffffffffffffff8ef3604401c",
    x"0802000000000000031ffffffffffffff6f669ea551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266df7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6431c",
    x"020900000000000000ae00000000000000fb3383691c",
    x"030b00000000000000aefffffffffffff50003e4991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd09c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f484d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd368f1c",
    x"070a00000000000000aefffffffffffff8ef36043d1c",
    x"080200000000000000aefffffffffffff6f669ea531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266df7b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6441c",
    x"020900000000000001a400000000000000fb3383631c",
    x"030b00000000000001a4fffffffffffff50003e49a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd09a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f48491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd36891c",
    x"070a00000000000001a4fffffffffffff8ef3604391c",
    x"080200000000000001a4fffffffffffff6f669ea501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266df771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe6451c",
    x"020900000000000001a600000000000000fb33835e1c",
    x"030b00000000000001a6fffffffffffff50003e49b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dd0981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f48451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd36831c",
    x"070a00000000000001a6fffffffffffff8ef3604361c",
    x"080200000000000001a6fffffffffffff6f669ea4e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6461c",
    x"0209000000000000015500000000000000fb3383581c",
    x"030b0000000000000155fffffffffffff50003e49c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd367c1c",
    x"070a0000000000000155fffffffffffff8ef3604321c",
    x"08020000000000000155fffffffffffff6f669ea4c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6471c",
    x"0209000000000000015500000000000000fb3383531c",
    x"030b0000000000000155fffffffffffff50003e49d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f483e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36761c",
    x"070a0000000000000155fffffffffffff8ef36042e1c",
    x"08020000000000000155fffffffffffff6f669ea491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6481c",
    x"0209000000000000015500000000000000fb33834d1c",
    x"030b0000000000000155fffffffffffff50003e49e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f483a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36701c",
    x"070a0000000000000155fffffffffffff8ef36042b1c",
    x"08020000000000000155fffffffffffff6f669ea471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6491c",
    x"0209000000000000015500000000000000fb3383471c",
    x"030b0000000000000155fffffffffffff50003e49f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd08e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd366a1c",
    x"070a0000000000000155fffffffffffff8ef3604271c",
    x"08020000000000000155fffffffffffff6f669ea451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe64a1c",
    x"0209000000000000015500000000000000fb3383421c",
    x"030b0000000000000155fffffffffffff50003e4a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd08c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48331c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36641c",
    x"070a0000000000000155fffffffffffff8ef3604241c",
    x"08020000000000000155fffffffffffff6f669ea421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df5e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe64b1c",
    x"0209000000000000015500000000000000fb33833c1c",
    x"030b0000000000000155fffffffffffff50003e4a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd08a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f482f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd365e1c",
    x"070a0000000000000155fffffffffffff8ef3604201c",
    x"08020000000000000155fffffffffffff6f669ea401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe64d1c",
    x"0209000000000000015500000000000000fb3383371c",
    x"030b0000000000000155fffffffffffff50003e4a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f482b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36581c",
    x"070a0000000000000155fffffffffffff8ef36041d1c",
    x"08020000000000000155fffffffffffff6f669ea3d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe64e1c",
    x"0209000000000000015500000000000000fb3383311c",
    x"030b0000000000000155fffffffffffff50003e4a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36521c",
    x"070a0000000000000155fffffffffffff8ef3604191c",
    x"08020000000000000155fffffffffffff6f669ea3b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe64f1c",
    x"0209000000000000015500000000000000fb33832b1c",
    x"030b0000000000000155fffffffffffff50003e4a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd364b1c",
    x"070a0000000000000155fffffffffffff8ef3604161c",
    x"08020000000000000155fffffffffffff6f669ea391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df4d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6501c",
    x"0209000000000000015500000000000000fb3383261c",
    x"030b0000000000000155fffffffffffff50003e4a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36451c",
    x"070a0000000000000155fffffffffffff8ef3604121c",
    x"08020000000000000155fffffffffffff6f669ea361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6511c",
    x"0209000000000000015500000000000000fb3383201c",
    x"030b0000000000000155fffffffffffff50003e4a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd07e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f481c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd363f1c",
    x"070a0000000000000155fffffffffffff8ef36040e1c",
    x"08020000000000000155fffffffffffff6f669ea341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6521c",
    x"0209000000000000015500000000000000fb33831b1c",
    x"030b0000000000000155fffffffffffff50003e4a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd07b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36391c",
    x"070a0000000000000155fffffffffffff8ef36040b1c",
    x"08020000000000000155fffffffffffff6f669ea321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6531c",
    x"0209000000000000015500000000000000fb3383151c",
    x"030b0000000000000155fffffffffffff50003e4a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36331c",
    x"070a0000000000000155fffffffffffff8ef3604071c",
    x"08020000000000000155fffffffffffff6f669ea2f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df3c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6541c",
    x"0209000000000000015500000000000000fb3383101c",
    x"030b0000000000000155fffffffffffff50003e4a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f48111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd362d1c",
    x"070a0000000000000155fffffffffffff8ef3604041c",
    x"08020000000000000155fffffffffffff6f669ea2d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266df381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe6551c",
    x"0209000000000000029500000000000000fb33830a1c",
    x"030b0000000000000295fffffffffffff50003e4aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd0741c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f480e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd36271c",
    x"070a0000000000000295fffffffffffff8ef3604001c",
    x"08020000000000000295fffffffffffff6f669ea2a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266df331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6561c",
    x"020900000000000002aa00000000000000fb3383041c",
    x"030b00000000000002aafffffffffffff50003e4ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0721c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f480a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd36201c",
    x"070a00000000000002aafffffffffffff8ef3603fd1c",
    x"080200000000000002aafffffffffffff6f669ea281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266df2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6571c",
    x"0209000000000000031f00000000000000fb3382ff1c",
    x"030b000000000000031ffffffffffffff50003e4ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd0701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f48061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd361a1c",
    x"070a000000000000031ffffffffffffff8ef3603f91c",
    x"0802000000000000031ffffffffffffff6f669ea261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266df2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6591c",
    x"020900000000000000ae00000000000000fb3382f91c",
    x"030b00000000000000aefffffffffffff50003e4ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd06d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f48021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd36141c",
    x"070a00000000000000aefffffffffffff8ef3603f51c",
    x"080200000000000000aefffffffffffff6f669ea231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266df271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe65a1c",
    x"020900000000000001a400000000000000fb3382f41c",
    x"030b00000000000001a4fffffffffffff50003e4ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd06b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f47ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd360e1c",
    x"070a00000000000001a4fffffffffffff8ef3603f21c",
    x"080200000000000001a4fffffffffffff6f669ea211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266df231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe65b1c",
    x"0209000000000000016600000000000000fb3382ee1c",
    x"030b0000000000000166fffffffffffff50003e4af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dd0681c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f47fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd36081c",
    x"070a0000000000000166fffffffffffff8ef3603ee1c",
    x"08020000000000000166fffffffffffff6f669ea1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe65c1c",
    x"0209000000000000015500000000000000fb3382e81c",
    x"030b0000000000000155fffffffffffff50003e4b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47f71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd36021c",
    x"070a0000000000000155fffffffffffff8ef3603eb1c",
    x"08020000000000000155fffffffffffff6f669ea1c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266df1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe65d1c",
    x"0209000000000000016500000000000000fb3382e31c",
    x"030b0000000000000165fffffffffffff50003e4b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dd0641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f47f31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd35fc1c",
    x"070a0000000000000165fffffffffffff8ef3603e71c",
    x"08020000000000000165fffffffffffff6f669ea1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe65e1c",
    x"0209000000000000015500000000000000fb3382dd1c",
    x"030b0000000000000155fffffffffffff50003e4b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35f61c",
    x"070a0000000000000155fffffffffffff8ef3603e41c",
    x"08020000000000000155fffffffffffff6f669ea171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe65f1c",
    x"0209000000000000015500000000000000fb3382d81c",
    x"030b0000000000000155fffffffffffff50003e4b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd05f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47ec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35ef1c",
    x"070a0000000000000155fffffffffffff8ef3603e01c",
    x"08020000000000000155fffffffffffff6f669ea151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df0e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6601c",
    x"0209000000000000015500000000000000fb3382d21c",
    x"030b0000000000000155fffffffffffff50003e4b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd05d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47e81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35e91c",
    x"070a0000000000000155fffffffffffff8ef3603dc1c",
    x"08020000000000000155fffffffffffff6f669ea131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6611c",
    x"0209000000000000015500000000000000fb3382cc1c",
    x"030b0000000000000155fffffffffffff50003e4b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd05a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47e51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35e31c",
    x"070a0000000000000155fffffffffffff8ef3603d91c",
    x"08020000000000000155fffffffffffff6f669ea101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6621c",
    x"0209000000000000015500000000000000fb3382c71c",
    x"030b0000000000000155fffffffffffff50003e4b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47e11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35dd1c",
    x"070a0000000000000155fffffffffffff8ef3603d51c",
    x"08020000000000000155fffffffffffff6f669ea0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266df011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6631c",
    x"0209000000000000015500000000000000fb3382c11c",
    x"030b0000000000000155fffffffffffff50003e4b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0561c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47dd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35d71c",
    x"070a0000000000000155fffffffffffff8ef3603d21c",
    x"08020000000000000155fffffffffffff6f669ea0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266defd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6651c",
    x"0209000000000000015500000000000000fb3382bc1c",
    x"030b0000000000000155fffffffffffff50003e4b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35d11c",
    x"070a0000000000000155fffffffffffff8ef3603ce1c",
    x"08020000000000000155fffffffffffff6f669ea091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266def91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6661c",
    x"0209000000000000015500000000000000fb3382b61c",
    x"030b0000000000000155fffffffffffff50003e4ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0511c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47d61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35cb1c",
    x"070a0000000000000155fffffffffffff8ef3603cb1c",
    x"08020000000000000155fffffffffffff6f669ea071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266def41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6671c",
    x"0209000000000000015500000000000000fb3382b11c",
    x"030b0000000000000155fffffffffffff50003e4bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd04e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47d21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35c51c",
    x"070a0000000000000155fffffffffffff8ef3603c71c",
    x"08020000000000000155fffffffffffff6f669ea041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266def01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6681c",
    x"0209000000000000015500000000000000fb3382ab1c",
    x"030b0000000000000155fffffffffffff50003e4bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd04c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35be1c",
    x"070a0000000000000155fffffffffffff8ef3603c31c",
    x"08020000000000000155fffffffffffff6f669ea021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266deec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6691c",
    x"0209000000000000015500000000000000fb3382a51c",
    x"030b0000000000000155fffffffffffff50003e4bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd04a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47cb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35b81c",
    x"070a0000000000000155fffffffffffff8ef3603c01c",
    x"08020000000000000155fffffffffffff6f669ea001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dee81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe66a1c",
    x"0209000000000000015500000000000000fb3382a01c",
    x"030b0000000000000155fffffffffffff50003e4be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47c71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35b21c",
    x"070a0000000000000155fffffffffffff8ef3603bc1c",
    x"08020000000000000155fffffffffffff6f669e9fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266dee41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe66b1c",
    x"0209000000000000025500000000000000fb33829a1c",
    x"030b0000000000000255fffffffffffff50003e4bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dd0451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f47c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd35ac1c",
    x"070a0000000000000255fffffffffffff8ef3603b91c",
    x"08020000000000000255fffffffffffff6f669e9fb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dedf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe66c1c",
    x"020900000000000002aa00000000000000fb3382951c",
    x"030b00000000000002aafffffffffffff50003e4c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35a61c",
    x"070a00000000000002aafffffffffffff8ef3603b51c",
    x"080200000000000002aafffffffffffff6f669e9f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dedb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe66d1c",
    x"0209000000000000031f00000000000000fb33828f1c",
    x"030b000000000000031ffffffffffffff50003e4c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd0401c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f47bc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd35a01c",
    x"070a000000000000031ffffffffffffff8ef3603b21c",
    x"0802000000000000031ffffffffffffff6f669e9f61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266ded71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe66e1c",
    x"020900000000000000ae00000000000000fb3382891c",
    x"030b00000000000000aefffffffffffff50003e4c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd03e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f47b81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd359a1c",
    x"070a00000000000000aefffffffffffff8ef3603ae1c",
    x"080200000000000000aefffffffffffff6f669e9f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ded31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe66f1c",
    x"020900000000000001a400000000000000fb3382841c",
    x"030b00000000000001a4fffffffffffff50003e4c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd03c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f47b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd35931c",
    x"070a00000000000001a4fffffffffffff8ef3603aa1c",
    x"080200000000000001a4fffffffffffff6f669e9f11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266decf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe6711c",
    x"0209000000000000026600000000000000fb33827e1c",
    x"030b0000000000000266fffffffffffff50003e4c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dd0391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f47b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000266ffffffffffffff04cd358d1c",
    x"070a0000000000000266fffffffffffff8ef3603a71c",
    x"08020000000000000266fffffffffffff6f669e9ef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266deca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6721c",
    x"020900000000000002aa00000000000000fb3382791c",
    x"030b00000000000002aafffffffffffff50003e4c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47ad1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35871c",
    x"070a00000000000002aafffffffffffff8ef3603a31c",
    x"080200000000000002aafffffffffffff6f669e9ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dec61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6731c",
    x"020900000000000002aa00000000000000fb3382731c",
    x"030b00000000000002aafffffffffffff50003e4c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47a91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35811c",
    x"070a00000000000002aafffffffffffff8ef3603a01c",
    x"080200000000000002aafffffffffffff6f669e9ea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dec21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6741c",
    x"020900000000000002aa00000000000000fb33826d1c",
    x"030b00000000000002aafffffffffffff50003e4c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd357b1c",
    x"070a00000000000002aafffffffffffff8ef36039c1c",
    x"080200000000000002aafffffffffffff6f669e9e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266debe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6751c",
    x"020900000000000002aa00000000000000fb3382681c",
    x"030b00000000000002aafffffffffffff50003e4c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0301c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47a21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35751c",
    x"070a00000000000002aafffffffffffff8ef3603991c",
    x"080200000000000002aafffffffffffff6f669e9e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266deba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6761c",
    x"020900000000000002aa00000000000000fb3382621c",
    x"030b00000000000002aafffffffffffff50003e4c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd02d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f479e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd356f1c",
    x"070a00000000000002aafffffffffffff8ef3603951c",
    x"080200000000000002aafffffffffffff6f669e9e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266deb51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6771c",
    x"020900000000000002aa00000000000000fb33825d1c",
    x"030b00000000000002aafffffffffffff50003e4ca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd02b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f479a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35681c",
    x"070a00000000000002aafffffffffffff8ef3603911c",
    x"080200000000000002aafffffffffffff6f669e9e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266deb11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6781c",
    x"020900000000000002aa00000000000000fb3382571c",
    x"030b00000000000002aafffffffffffff50003e4cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0291c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35621c",
    x"070a00000000000002aafffffffffffff8ef36038e1c",
    x"080200000000000002aafffffffffffff6f669e9de1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dead1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6791c",
    x"020900000000000002aa00000000000000fb3382511c",
    x"030b00000000000002aafffffffffffff50003e4cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd355c1c",
    x"070a00000000000002aafffffffffffff8ef36038a1c",
    x"080200000000000002aafffffffffffff6f669e9dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dea91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe67a1c",
    x"020900000000000002aa00000000000000fb33824c1c",
    x"030b00000000000002aafffffffffffff50003e4cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f478f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35561c",
    x"070a00000000000002aafffffffffffff8ef3603871c",
    x"080200000000000002aafffffffffffff6f669e9da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dea51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe67b1c",
    x"020900000000000002aa00000000000000fb3382461c",
    x"030b00000000000002aafffffffffffff50003e4cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f478b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35501c",
    x"070a00000000000002aafffffffffffff8ef3603831c",
    x"080200000000000002aafffffffffffff6f669e9d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dea01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe67d1c",
    x"020900000000000002aa00000000000000fb3382411c",
    x"030b00000000000002aafffffffffffff50003e4d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd01f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd354a1c",
    x"070a00000000000002aafffffffffffff8ef3603801c",
    x"080200000000000002aafffffffffffff6f669e9d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266de9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe67e1c",
    x"020900000000000002aa00000000000000fb33823b1c",
    x"030b00000000000002aafffffffffffff50003e4d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd01d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35441c",
    x"070a00000000000002aafffffffffffff8ef36037c1c",
    x"080200000000000002aafffffffffffff6f669e9d31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266de981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe67f1c",
    x"020900000000000002aa00000000000000fb3382361c",
    x"030b00000000000002aafffffffffffff50003e4d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd01a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd353e1c",
    x"070a00000000000002aafffffffffffff8ef3603791c",
    x"080200000000000002aafffffffffffff6f669e9d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266de941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6801c",
    x"020900000000000002aa00000000000000fb3382301c",
    x"030b00000000000002aafffffffffffff50003e4d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f477c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35371c",
    x"070a00000000000002aafffffffffffff8ef3603751c",
    x"080200000000000002aafffffffffffff6f669e9ce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266de901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6811c",
    x"020900000000000002aa00000000000000fb33822a1c",
    x"030b00000000000002aafffffffffffff50003e4d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd35311c",
    x"070a00000000000002aafffffffffffff8ef3603711c",
    x"080200000000000002aafffffffffffff6f669e9cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266de8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6821c",
    x"020900000000000002aa00000000000000fb3382251c",
    x"030b00000000000002aafffffffffffff50003e4d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dd0131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd352b1c",
    x"070a00000000000002aafffffffffffff8ef36036e1c",
    x"080200000000000002aafffffffffffff6f669e9c91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266de871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6831c",
    x"0209000000000000031f00000000000000fb33821f1c",
    x"030b000000000000031ffffffffffffff50003e4d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dd0111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f47711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd35251c",
    x"070a000000000000031ffffffffffffff8ef36036a1c",
    x"0802000000000000031ffffffffffffff6f669e9c71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266de831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6841c",
    x"020900000000000000ae00000000000000fb33821a1c",
    x"030b00000000000000aefffffffffffff50003e4d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dd00f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f476e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd351f1c",
    x"070a00000000000000aefffffffffffff8ef3603671c",
    x"080200000000000000aefffffffffffff6f669e9c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266de7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6851c",
    x"020900000000000001a400000000000000fb3382141c",
    x"030b00000000000001a4fffffffffffff50003e4d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dd00c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f476a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd35191c",
    x"070a00000000000001a4fffffffffffff8ef3603631c",
    x"080200000000000001a4fffffffffffff6f669e9c21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266de7b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbe6861c",
    x"020900000000000001aa00000000000000fb33820e1c",
    x"030b00000000000001aafffffffffffff50003e4d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dd00a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f47661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd35131c",
    x"070a00000000000001aafffffffffffff8ef3603601c",
    x"080200000000000001aafffffffffffff6f669e9c01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266de761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe6871c",
    x"0209000000000000029500000000000000fb3382091c",
    x"030b0000000000000295fffffffffffff50003e4da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dd0071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f47621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd350c1c",
    x"070a0000000000000295fffffffffffff8ef36035c1c",
    x"08020000000000000295fffffffffffff6f669e9bd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266de721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe6891c",
    x"0209000000000000015a00000000000000fb3382031c",
    x"030b000000000000015afffffffffffff50003e4db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dd0051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f475f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd35061c",
    x"070a000000000000015afffffffffffff8ef3603581c",
    x"0802000000000000015afffffffffffff6f669e9bb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266de6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe68a1c",
    x"0209000000000000015500000000000000fb3381fe1c",
    x"030b0000000000000155fffffffffffff50003e4dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dd0031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f475b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd35001c",
    x"070a0000000000000155fffffffffffff8ef3603551c",
    x"08020000000000000155fffffffffffff6f669e9b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266de6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe68b1c",
    x"0209000000000000015600000000000000fb3381f81c",
    x"030b00000000000002aafffffffffffff50003e4dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dd0001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd34fa1c",
    x"070a00000000000002aafffffffffffff8ef3603511c",
    x"08020000000000000156fffffffffffff6f669e9b61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266de661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe68c1c",
    x"0209000000000000016500000000000000fb3381f21c",
    x"030b000000000000019afffffffffffff50003e4de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcffe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a90000000000000b072f47531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd34f41c",
    x"070a00000000000001aafffffffffffff8ef36034e1c",
    x"08020000000000000156fffffffffffff6f669e9b41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266de611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe68d1c",
    x"020900000000000002a500000000000000fb3381ed1c",
    x"030b000000000000019afffffffffffff50003e4df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcffc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd34ee1c",
    x"070a0000000000000165fffffffffffff8ef36034a1c",
    x"08020000000000000265fffffffffffff6f669e9b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266de5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe68e1c",
    x"0209000000000000026600000000000000fb3381e71c",
    x"030b0000000000000299fffffffffffff50003e4e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dcff91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f474c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd34e81c",
    x"070a0000000000000256fffffffffffff8ef3603471c",
    x"08020000000000000195fffffffffffff6f669e9af1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266de591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe68f1c",
    x"0209000000000000029900000000000000fb3381e21c",
    x"030b0000000000000259fffffffffffff50003e4e11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcff71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f47481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd34e21c",
    x"070a0000000000000266fffffffffffff8ef3603431c",
    x"080200000000000001a5fffffffffffff6f669e9ad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266de551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6901c",
    x"020900000000000002aa00000000000000fb3381dc1c",
    x"030b00000000000002a5fffffffffffff50003e4e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dcff41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f47451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd34db1c",
    x"070a0000000000000295fffffffffffff8ef36033f1c",
    x"080200000000000001a5fffffffffffff6f669e9aa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266de511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe6911c",
    x"020900000000000002a500000000000000fb3381d61c",
    x"030b000000000000016afffffffffffff50003e4e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcff21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f47411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd34d51c",
    x"070a0000000000000255fffffffffffff8ef36033c1c",
    x"08020000000000000169fffffffffffff6f669e9a81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266de4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe6921c",
    x"0209000000000000025600000000000000fb3381d11c",
    x"030b0000000000000166fffffffffffff50003e4e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcff01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f473d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd34cf1c",
    x"070a000000000000029afffffffffffff8ef3603381c",
    x"08020000000000000295fffffffffffff6f669e9a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000269ffffffffffffff0266de481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbe6931c",
    x"0209000000000000015500000000000000fb3381cb1c",
    x"030b0000000000000296fffffffffffff50003e4e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dcfed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f47391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd34c91c",
    x"070a0000000000000156fffffffffffff8ef3603351c",
    x"08020000000000000266fffffffffffff6f669e9a31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266de441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe6951c",
    x"0209000000000000016500000000000000fb3381c61c",
    x"030b0000000000000265fffffffffffff50003e4e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dcfeb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f47361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000265ffffffffffffff04cd34c31c",
    x"070a0000000000000295fffffffffffff8ef3603311c",
    x"0802000000000000029afffffffffffff6f669e9a11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266de401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a90000000000000b0bfbe6961c",
    x"0209000000000000015900000000000000fb3381c01c",
    x"030b00000000000002a5fffffffffffff50003e4e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dcfe91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f47321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd34bd1c",
    x"070a00000000000001a5fffffffffffff8ef36032d1c",
    x"080200000000000001a5fffffffffffff6f669e99e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266de3c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a90000000000000b0bfbe6971c",
    x"0209000000000000029500000000000000fb3381bb1c",
    x"030b000000000000025afffffffffffff50003e4e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dcfe61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f472e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd34b71c",
    x"070a0000000000000166fffffffffffff8ef36032a1c",
    x"08020000000000000196fffffffffffff6f669e99c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266de371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6981c",
    x"020900000000000002a500000000000000fb3381b51c",
    x"030b000000000000015afffffffffffff50003e4e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcfe41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f472b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd34b01c",
    x"070a000000000000015afffffffffffff8ef3603261c",
    x"08020000000000000296fffffffffffff6f669e99a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266de331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6991c",
    x"0209000000000000031f00000000000000fb3381af1c",
    x"030b000000000000031ffffffffffffff50003e4ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcfe21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f47271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd34aa1c",
    x"070a000000000000031ffffffffffffff8ef3603231c",
    x"0802000000000000031ffffffffffffff6f669e9971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266de2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe69a1c",
    x"020900000000000000ae00000000000000fb3381aa1c",
    x"030b00000000000000aefffffffffffff50003e4eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcfdf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f47231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd34a41c",
    x"070a00000000000000aefffffffffffff8ef36031f1c",
    x"080200000000000000aefffffffffffff6f669e9951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266de2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe69b1c",
    x"020900000000000001a400000000000000fb3381a41c",
    x"030b00000000000001a4fffffffffffff50003e4ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcfdd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f471f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd349e1c",
    x"070a00000000000001a4fffffffffffff8ef36031c1c",
    x"080200000000000001a4fffffffffffff6f669e9921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266de271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe69c1c",
    x"0209000000000000016a00000000000000fb33819f1c",
    x"030b000000000000016afffffffffffff50003e4ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcfda1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f471c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd34981c",
    x"070a000000000000016afffffffffffff8ef3603181c",
    x"0802000000000000016afffffffffffff6f669e9901c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266de221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe69d1c",
    x"0209000000000000015500000000000000fb3381991c",
    x"030b0000000000000155fffffffffffff50003e4ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcfd81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f47181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd34921c",
    x"070a0000000000000155fffffffffffff8ef3603141c",
    x"08020000000000000155fffffffffffff6f669e98e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266de1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe69e1c",
    x"0209000000000000019500000000000000fb3381931c",
    x"030b0000000000000195fffffffffffff50003e4ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dcfd61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f47141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd348c1c",
    x"070a0000000000000195fffffffffffff8ef3603111c",
    x"080200000000000002a5fffffffffffff6f669e98b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266de1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6a01c",
    x"020900000000000002aa00000000000000fb33818e1c",
    x"030b00000000000002aafffffffffffff50003e4f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcfd31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f47111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd34851c",
    x"070a00000000000002aafffffffffffff8ef36030d1c",
    x"08020000000000000155fffffffffffff6f669e9891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266de161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe6a11c",
    x"0209000000000000029600000000000000fb3381881c",
    x"030b00000000000001aafffffffffffff50003e4f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcfd11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f470d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd347f1c",
    x"070a0000000000000256fffffffffffff8ef36030a1c",
    x"08020000000000000155fffffffffffff6f669e9871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266de121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe6a21c",
    x"0209000000000000026500000000000000fb3381831c",
    x"030b00000000000002a9fffffffffffff50003e4f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dcfcf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f47091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd34791c",
    x"070a000000000000029afffffffffffff8ef3603061c",
    x"08020000000000000159fffffffffffff6f669e9841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266de0d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe6a31c",
    x"0209000000000000029600000000000000fb33817d1c",
    x"030b000000000000016afffffffffffff50003e4f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dcfcc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f47051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd34731c",
    x"070a0000000000000159fffffffffffff8ef3603031c",
    x"0802000000000000015afffffffffffff6f669e9821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266de091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6a41c",
    x"0209000000000000016900000000000000fb3381771c",
    x"030b0000000000000295fffffffffffff50003e4f51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcfca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f47021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd346d1c",
    x"070a0000000000000196fffffffffffff8ef3602ff1c",
    x"08020000000000000299fffffffffffff6f669e97f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266de051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe6a51c",
    x"020900000000000002a500000000000000fb3381721c",
    x"030b0000000000000156fffffffffffff50003e4f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dcfc71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f46fe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd34671c",
    x"070a00000000000002a6fffffffffffff8ef3602fb1c",
    x"080200000000000001a5fffffffffffff6f669e97d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266de011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe6a61c",
    x"0209000000000000025500000000000000fb33816c1c",
    x"030b000000000000016afffffffffffff50003e4f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcfc51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f46fa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd34611c",
    x"070a0000000000000295fffffffffffff8ef3602f81c",
    x"0802000000000000026afffffffffffff6f669e97b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266ddfd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe6a71c",
    x"0209000000000000029a00000000000000fb3381671c",
    x"030b0000000000000269fffffffffffff50003e4f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dcfc31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f46f71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd345b1c",
    x"070a0000000000000196fffffffffffff8ef3602f41c",
    x"08020000000000000165fffffffffffff6f669e9781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ddf81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe6a81c",
    x"020900000000000001a600000000000000fb3381611c",
    x"030b000000000000019afffffffffffff50003e4f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcfc01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f46f31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd34541c",
    x"070a000000000000026afffffffffffff8ef3602f11c",
    x"0802000000000000019afffffffffffff6f669e9761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266ddf41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbe6a91c",
    x"0209000000000000025a00000000000000fb33815b1c",
    x"030b00000000000002a9fffffffffffff50003e4fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcfbe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f46ef1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd344e1c",
    x"070a00000000000002a6fffffffffffff8ef3602ed1c",
    x"08020000000000000295fffffffffffff6f669e9741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266ddf01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe6aa1c",
    x"0209000000000000029600000000000000fb3381561c",
    x"030b000000000000025afffffffffffff50003e4fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dcfbc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f46eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd34481c",
    x"070a000000000000019afffffffffffff8ef3602ea1c",
    x"0802000000000000029afffffffffffff6f669e9711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266ddec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe6ac1c",
    x"0209000000000000019900000000000000fb3381501c",
    x"030b0000000000000156fffffffffffff50003e4fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcfb91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f46e81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd34421c",
    x"070a0000000000000166fffffffffffff8ef3602e61c",
    x"080200000000000001a9fffffffffffff6f669e96f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266dde81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe6ad1c",
    x"0209000000000000015600000000000000fb33814b1c",
    x"030b0000000000000169fffffffffffff50003e4fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcfb71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f46e41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd343c1c",
    x"070a0000000000000159fffffffffffff8ef3602e21c",
    x"08020000000000000255fffffffffffff6f669e96c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266dde31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6ae1c",
    x"0209000000000000029a00000000000000fb3381451c",
    x"030b00000000000002a9fffffffffffff50003e4fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcfb41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46e01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd34361c",
    x"070a0000000000000159fffffffffffff8ef3602df1c",
    x"08020000000000000299fffffffffffff6f669e96a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dddf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6af1c",
    x"0209000000000000031f00000000000000fb3381401c",
    x"030b000000000000031ffffffffffffff50003e4ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcfb21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f46dd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd34301c",
    x"070a000000000000031ffffffffffffff8ef3602db1c",
    x"0802000000000000031ffffffffffffff6f669e9681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dddb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6b01c",
    x"020900000000000000ae00000000000000fb33813a1c",
    x"030b00000000000000aefffffffffffff50003e5001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcfb01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f46d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd34291c",
    x"070a00000000000000aefffffffffffff8ef3602d81c",
    x"080200000000000000aefffffffffffff6f669e9651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ddd71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6b11c",
    x"020900000000000001a400000000000000fb3381341c",
    x"030b00000000000001a4fffffffffffff50003e5011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcfad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f46d51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd34231c",
    x"070a00000000000001a4fffffffffffff8ef3602d41c",
    x"080200000000000001a4fffffffffffff6f669e9631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266ddd31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe6b21c",
    x"0209000000000000026a00000000000000fb33812f1c",
    x"030b000000000000026afffffffffffff50003e5021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dcfab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f46d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026affffffffffffff04cd341d1c",
    x"070a000000000000026afffffffffffff8ef3602d11c",
    x"0802000000000000026afffffffffffff6f669e9611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ddce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6b31c",
    x"0209000000000000015500000000000000fb3381291c",
    x"030b0000000000000155fffffffffffff50003e5031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcfa91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f46ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd34171c",
    x"070a00000000000002a9fffffffffffff8ef3602cd1c",
    x"08020000000000000155fffffffffffff6f669e95e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ddca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6b41c",
    x"0209000000000000015500000000000000fb3381241c",
    x"030b0000000000000155fffffffffffff50003e5041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcfa61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f46ca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd34111c",
    x"070a00000000000001aafffffffffffff8ef3602c91c",
    x"08020000000000000155fffffffffffff6f669e95c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266ddc61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe6b51c",
    x"0209000000000000015600000000000000fb33811e1c",
    x"030b0000000000000155fffffffffffff50003e5051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dcfa41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f46c61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd340b1c",
    x"070a00000000000002aafffffffffffff8ef3602c61c",
    x"08020000000000000155fffffffffffff6f669e9591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ddc21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe6b61c",
    x"0209000000000000025500000000000000fb3381181c",
    x"030b0000000000000195fffffffffffff50003e5061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcfa11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f46c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd34051c",
    x"070a000000000000026afffffffffffff8ef3602c21c",
    x"08020000000000000195fffffffffffff6f669e9571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266ddbe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe6b81c",
    x"0209000000000000016500000000000000fb3381131c",
    x"030b00000000000002a9fffffffffffff50003e5071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dcf9f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000259ffffffffffffff04cd33ff1c",
    x"070a0000000000000256fffffffffffff8ef3602bf1c",
    x"08020000000000000299fffffffffffff6f669e9551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266ddb91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe6b91c",
    x"0209000000000000019900000000000000fb33810d1c",
    x"030b0000000000000195fffffffffffff50003e5081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dcf9d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f46bb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd33f81c",
    x"070a0000000000000266fffffffffffff8ef3602bb1c",
    x"080200000000000002a6fffffffffffff6f669e9521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266ddb51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe6ba1c",
    x"0209000000000000016500000000000000fb3381081c",
    x"030b0000000000000166fffffffffffff50003e5091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dcf9a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f46b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd33f21c",
    x"070a0000000000000156fffffffffffff8ef3602b81c",
    x"0802000000000000025afffffffffffff6f669e9501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266ddb11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe6bb1c",
    x"0209000000000000019500000000000000fb3381021c",
    x"030b0000000000000265fffffffffffff50003e50a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dcf981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f46b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd33ec1c",
    x"070a000000000000025afffffffffffff8ef3602b41c",
    x"0802000000000000016afffffffffffff6f669e94e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ddad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe6bc1c",
    x"0209000000000000026a00000000000000fb3380fc1c",
    x"030b00000000000002aafffffffffffff50003e50b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f46b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd33e61c",
    x"070a0000000000000195fffffffffffff8ef3602b01c",
    x"08020000000000000195fffffffffffff6f669e94b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266dda91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe6bd1c",
    x"0209000000000000025600000000000000fb3380f71c",
    x"030b00000000000002a5fffffffffffff50003e50c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dcf931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f46ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd33e01c",
    x"070a00000000000002a5fffffffffffff8ef3602ad1c",
    x"08020000000000000295fffffffffffff6f669e9491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266dda41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe6be1c",
    x"020900000000000001a900000000000000fb3380f11c",
    x"030b0000000000000155fffffffffffff50003e50d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dcf911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f46a91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd33da1c",
    x"070a0000000000000256fffffffffffff8ef3602a91c",
    x"08020000000000000199fffffffffffff6f669e9461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266dda01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe6bf1c",
    x"0209000000000000029500000000000000fb3380ec1c",
    x"030b0000000000000299fffffffffffff50003e50e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf8f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f46a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd33d41c",
    x"070a0000000000000266fffffffffffff8ef3602a61c",
    x"08020000000000000166fffffffffffff6f669e9441c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266dd9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe6c01c",
    x"0209000000000000016900000000000000fb3380e61c",
    x"030b000000000000016afffffffffffff50003e50f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dcf8c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f46a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd33cd1c",
    x"070a0000000000000256fffffffffffff8ef3602a21c",
    x"08020000000000000199fffffffffffff6f669e9421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266dd981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe6c11c",
    x"0209000000000000026a00000000000000fb3380e01c",
    x"030b000000000000016afffffffffffff50003e5101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dcf8a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f469d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd33c71c",
    x"070a00000000000001a5fffffffffffff8ef36029e1c",
    x"08020000000000000266fffffffffffff6f669e93f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266dd941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe6c31c",
    x"020900000000000001a900000000000000fb3380db1c",
    x"030b000000000000026afffffffffffff50003e5111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dcf871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f469a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd33c11c",
    x"070a0000000000000166fffffffffffff8ef36029b1c",
    x"08020000000000000296fffffffffffff6f669e93d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266dd8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe6c41c",
    x"020900000000000002a600000000000000fb3380d51c",
    x"030b000000000000015afffffffffffff50003e5121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dcf851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f46961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd33bb1c",
    x"070a0000000000000295fffffffffffff8ef3602971c",
    x"080200000000000002a5fffffffffffff6f669e93b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dd8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6c51c",
    x"0209000000000000031f00000000000000fb3380d01c",
    x"030b000000000000031ffffffffffffff50003e5131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcf831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f46921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd33b51c",
    x"070a000000000000031ffffffffffffff8ef3602941c",
    x"0802000000000000031ffffffffffffff6f669e9381c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dd871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6c61c",
    x"020900000000000000ae00000000000000fb3380ca1c",
    x"030b00000000000000aefffffffffffff50003e5141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcf801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f468f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd33af1c",
    x"070a00000000000000aefffffffffffff8ef3602901c",
    x"080200000000000000aefffffffffffff6f669e9361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dd831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6c71c",
    x"020900000000000001a400000000000000fb3380c51c",
    x"030b00000000000001a4fffffffffffff50003e5161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcf7e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f468b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd33a91c",
    x"070a00000000000001a4fffffffffffff8ef36028d1c",
    x"080200000000000001a4fffffffffffff6f669e9331c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266dd7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe6c81c",
    x"0209000000000000015a00000000000000fb3380bf1c",
    x"030b000000000000015afffffffffffff50003e5171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dcf7c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f46871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd33a21c",
    x"070a000000000000015afffffffffffff8ef3602891c",
    x"0802000000000000015afffffffffffff6f669e9311c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd7a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6c91c",
    x"020900000000000001aa00000000000000fb3380b91c",
    x"030b0000000000000255fffffffffffff50003e5181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46831c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd339c1c",
    x"070a0000000000000155fffffffffffff8ef3602851c",
    x"08020000000000000155fffffffffffff6f669e92f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266dd761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe6ca1c",
    x"0209000000000000016900000000000000fb3380b41c",
    x"030b0000000000000269fffffffffffff50003e5191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dcf771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f46801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd33961c",
    x"070a00000000000002a6fffffffffffff8ef3602821c",
    x"080200000000000001a5fffffffffffff6f669e92c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266dd721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe6cb1c",
    x"020900000000000001a600000000000000fb3380ae1c",
    x"030b0000000000000296fffffffffffff50003e51a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dcf741c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f467c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd33901c",
    x"070a000000000000029afffffffffffff8ef36027e1c",
    x"08020000000000000196fffffffffffff6f669e92a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266dd6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe6cc1c",
    x"0209000000000000026900000000000000fb3380a91c",
    x"030b0000000000000255fffffffffffff50003e51b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dcf721c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f46781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000199ffffffffffffff04cd338a1c",
    x"070a0000000000000265fffffffffffff8ef36027b1c",
    x"08020000000000000256fffffffffffff6f669e9281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe6cd1c",
    x"0209000000000000015600000000000000fb3380a31c",
    x"030b0000000000000155fffffffffffff50003e51c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f46751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd33841c",
    x"070a00000000000002aafffffffffffff8ef3602771c",
    x"08020000000000000155fffffffffffff6f669e9251c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266dd651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbe6cf1c",
    x"0209000000000000025500000000000000fb33809d1c",
    x"030b0000000000000255fffffffffffff50003e51d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcf6d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f46711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd337e1c",
    x"070a00000000000001aafffffffffffff8ef3602741c",
    x"08020000000000000255fffffffffffff6f669e9231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dd611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6d01c",
    x"020900000000000002aa00000000000000fb3380981c",
    x"030b00000000000002aafffffffffffff50003e51e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf6b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f466d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33781c",
    x"070a0000000000000155fffffffffffff8ef3602701c",
    x"080200000000000002aafffffffffffff6f669e9201c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dd5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6d11c",
    x"020900000000000002aa00000000000000fb3380921c",
    x"030b00000000000002aafffffffffffff50003e51f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33711c",
    x"070a0000000000000155fffffffffffff8ef36026c1c",
    x"080200000000000002aafffffffffffff6f669e91e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dd591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6d21c",
    x"020900000000000002aa00000000000000fb33808d1c",
    x"030b00000000000002aafffffffffffff50003e5201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd336b1c",
    x"070a0000000000000155fffffffffffff8ef3602691c",
    x"080200000000000002aafffffffffffff6f669e91c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266dd551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbe6d31c",
    x"020900000000000001a600000000000000fb3380871c",
    x"030b00000000000001a6fffffffffffff50003e5211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000259fffffffffffff4099dcf641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f46621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd33651c",
    x"070a0000000000000259fffffffffffff8ef3602651c",
    x"080200000000000001a6fffffffffffff6f669e9191c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dd501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6d41c",
    x"020900000000000002aa00000000000000fb3380811c",
    x"030b00000000000002aafffffffffffff50003e5221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f465e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd335f1c",
    x"070a0000000000000155fffffffffffff8ef3602621c",
    x"080200000000000002aafffffffffffff6f669e9171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dd4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6d51c",
    x"020900000000000002aa00000000000000fb33807c1c",
    x"030b00000000000002aafffffffffffff50003e5231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf5f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f465b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33591c",
    x"070a0000000000000155fffffffffffff8ef36025e1c",
    x"080200000000000002aafffffffffffff6f669e9141c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266dd481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe6d61c",
    x"020900000000000002a600000000000000fb3380761c",
    x"030b00000000000002a6fffffffffffff50003e5241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcf5d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f46571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd33531c",
    x"070a0000000000000159fffffffffffff8ef36025a1c",
    x"080200000000000002a6fffffffffffff6f669e9121c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266dd441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a50000000000000b0bfbe6d71c",
    x"0209000000000000029500000000000000fb3380711c",
    x"030b00000000000002aafffffffffffff50003e5251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dcf5a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f46531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd334d1c",
    x"070a000000000000019afffffffffffff8ef3602571c",
    x"080200000000000002a5fffffffffffff6f669e9101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266dd401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe6d81c",
    x"0209000000000000015a00000000000000fb33806b1c",
    x"030b000000000000015afffffffffffff50003e5261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dcf581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f464f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd33461c",
    x"070a0000000000000255fffffffffffff8ef3602531c",
    x"0802000000000000019afffffffffffff6f669e90d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266dd3b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe6d91c",
    x"0209000000000000015a00000000000000fb3380651c",
    x"030b000000000000015afffffffffffff50003e5271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dcf561c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f464c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd33401c",
    x"070a00000000000002a5fffffffffffff8ef3602501c",
    x"0802000000000000015afffffffffffff6f669e90b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dd371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6db1c",
    x"0209000000000000031f00000000000000fb3380601c",
    x"030b000000000000031ffffffffffffff50003e5281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcf531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f46481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd333a1c",
    x"070a000000000000031ffffffffffffff8ef36024c1c",
    x"0802000000000000031ffffffffffffff6f669e9091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dd331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6dc1c",
    x"020900000000000000ae00000000000000fb33805a1c",
    x"030b00000000000000aefffffffffffff50003e5291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcf511c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f46441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd33341c",
    x"070a00000000000000aefffffffffffff8ef3602491c",
    x"080200000000000000aefffffffffffff6f669e9061c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dd2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6dd1c",
    x"020900000000000001a400000000000000fb3380551c",
    x"030b00000000000001a4fffffffffffff50003e52a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcf4e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f46411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd332e1c",
    x"070a00000000000001a4fffffffffffff8ef3602451c",
    x"080200000000000001a4fffffffffffff6f669e9041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266dd2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe6de1c",
    x"0209000000000000025a00000000000000fb33804f1c",
    x"030b000000000000025afffffffffffff50003e52b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dcf4c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f463d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd33281c",
    x"070a000000000000025afffffffffffff8ef3602411c",
    x"0802000000000000025afffffffffffff6f669e9011c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6df1c",
    x"020900000000000002aa00000000000000fb33804a1c",
    x"030b00000000000002aafffffffffffff50003e52c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf4a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f46391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33221c",
    x"070a00000000000002aafffffffffffff8ef36023e1c",
    x"080200000000000002aafffffffffffff6f669e8ff1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266dd221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe6e01c",
    x"0209000000000000029a00000000000000fb3380441c",
    x"030b000000000000029afffffffffffff50003e52d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcf471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f46351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd331b1c",
    x"070a000000000000029afffffffffffff8ef36023a1c",
    x"0802000000000000029afffffffffffff6f669e8fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e11c",
    x"020900000000000002aa00000000000000fb33803e1c",
    x"030b00000000000002aafffffffffffff50003e52e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f46321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33151c",
    x"070a00000000000002aafffffffffffff8ef3602371c",
    x"080200000000000002aafffffffffffff6f669e8fa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e21c",
    x"020900000000000002aa00000000000000fb3380391c",
    x"030b00000000000002aafffffffffffff50003e52f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f462e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd330f1c",
    x"070a00000000000002aafffffffffffff8ef3602331c",
    x"080200000000000002aafffffffffffff6f669e8f81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e31c",
    x"020900000000000002aa00000000000000fb3380331c",
    x"030b00000000000002aafffffffffffff50003e5301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf401c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f462a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33091c",
    x"070a00000000000002aafffffffffffff8ef3602301c",
    x"080200000000000002aafffffffffffff6f669e8f61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e41c",
    x"020900000000000002aa00000000000000fb33802e1c",
    x"030b00000000000002aafffffffffffff50003e5311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf3e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f46271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd33031c",
    x"070a00000000000002aafffffffffffff8ef36022c1c",
    x"080200000000000002aafffffffffffff6f669e8f31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd0d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e61c",
    x"020900000000000002aa00000000000000fb3380281c",
    x"030b00000000000002aafffffffffffff50003e5321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf3b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f46231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32fd1c",
    x"070a00000000000002aafffffffffffff8ef3602281c",
    x"080200000000000002aafffffffffffff6f669e8f11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e71c",
    x"020900000000000002aa00000000000000fb3380221c",
    x"030b00000000000002aafffffffffffff50003e5331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f461f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32f71c",
    x"070a00000000000002aafffffffffffff8ef3602251c",
    x"080200000000000002aafffffffffffff6f669e8ee1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dd051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6e81c",
    x"020900000000000002aa00000000000000fb33801d1c",
    x"030b00000000000002aafffffffffffff50003e5341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f461b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32f01c",
    x"070a00000000000002aafffffffffffff8ef3602211c",
    x"080200000000000002aafffffffffffff6f669e8ec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266dd011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe6e91c",
    x"0209000000000000016600000000000000fb3380171c",
    x"030b0000000000000166fffffffffffff50003e5351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dcf341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f46181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd32ea1c",
    x"070a0000000000000166fffffffffffff8ef36021e1c",
    x"08020000000000000166fffffffffffff6f669e8ea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dcfc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6ea1c",
    x"0209000000000000015500000000000000fb3380121c",
    x"030b0000000000000155fffffffffffff50003e5361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32e41c",
    x"070a0000000000000155fffffffffffff8ef36021a1c",
    x"08020000000000000155fffffffffffff6f669e8e71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dcf81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6eb1c",
    x"0209000000000000015500000000000000fb33800c1c",
    x"030b0000000000000155fffffffffffff50003e5371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf2f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46101c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32de1c",
    x"070a0000000000000155fffffffffffff8ef3602161c",
    x"08020000000000000155fffffffffffff6f669e8e51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dcf41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6ec1c",
    x"0209000000000000015500000000000000fb3380061c",
    x"030b0000000000000155fffffffffffff50003e5381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf2d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f460d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32d81c",
    x"070a0000000000000155fffffffffffff8ef3602131c",
    x"08020000000000000155fffffffffffff6f669e8e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dcf01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6ed1c",
    x"0209000000000000015500000000000000fb3380011c",
    x"030b0000000000000155fffffffffffff50003e5391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf2b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32d21c",
    x"070a0000000000000155fffffffffffff8ef36020f1c",
    x"08020000000000000155fffffffffffff6f669e8e01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dcec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe6ee1c",
    x"0209000000000000015500000000000000fb337ffb1c",
    x"030b0000000000000155fffffffffffff50003e53a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcf281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f46051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32cc1c",
    x"070a0000000000000155fffffffffffff8ef36020c1c",
    x"08020000000000000155fffffffffffff6f669e8de1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266dce71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe6ef1c",
    x"0209000000000000015900000000000000fb337ff61c",
    x"030b0000000000000159fffffffffffff50003e53b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcf261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f46011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd32c61c",
    x"070a0000000000000159fffffffffffff8ef3602081c",
    x"08020000000000000159fffffffffffff6f669e8db1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dce31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe6f01c",
    x"0209000000000000031f00000000000000fb337ff01c",
    x"030b000000000000031ffffffffffffff50003e53c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcf241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f45fe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd32bf1c",
    x"070a000000000000031ffffffffffffff8ef3602051c",
    x"0802000000000000031ffffffffffffff6f669e8d91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dcdf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe6f21c",
    x"020900000000000000ae00000000000000fb337fea1c",
    x"030b00000000000000aefffffffffffff50003e53d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcf211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f45fa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd32b91c",
    x"070a00000000000000aefffffffffffff8ef3602011c",
    x"080200000000000000aefffffffffffff6f669e8d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dcdb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe6f31c",
    x"020900000000000001a400000000000000fb337fe51c",
    x"030b00000000000001a4fffffffffffff50003e53e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcf1f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f45f61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd32b31c",
    x"070a00000000000001a4fffffffffffff8ef3601fd1c",
    x"080200000000000001a4fffffffffffff6f669e8d41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266dcd71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe6f41c",
    x"0209000000000000029a00000000000000fb337fdf1c",
    x"030b000000000000029afffffffffffff50003e53f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcf1c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f45f31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd32ad1c",
    x"070a000000000000029afffffffffffff8ef3601fa1c",
    x"0802000000000000029afffffffffffff6f669e8d21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266dcd21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe6f51c",
    x"0209000000000000016a00000000000000fb337fda1c",
    x"030b000000000000016afffffffffffff50003e5411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcf1a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f45ef1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd32a71c",
    x"070a000000000000016afffffffffffff8ef3601f61c",
    x"0802000000000000016afffffffffffff6f669e8d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6f61c",
    x"020900000000000002aa00000000000000fb337fd41c",
    x"030b00000000000002aafffffffffffff50003e5421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32a11c",
    x"070a00000000000002aafffffffffffff8ef3601f31c",
    x"080200000000000002aafffffffffffff6f669e8cd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6f71c",
    x"020900000000000002aa00000000000000fb337fce1c",
    x"030b00000000000002aafffffffffffff50003e5431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45e71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd329b1c",
    x"070a00000000000002aafffffffffffff8ef3601ef1c",
    x"080200000000000002aafffffffffffff6f669e8cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcc61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6f81c",
    x"020900000000000002aa00000000000000fb337fc91c",
    x"030b00000000000002aafffffffffffff50003e5441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45e41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32941c",
    x"070a00000000000002aafffffffffffff8ef3601eb1c",
    x"080200000000000002aafffffffffffff6f669e8c81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcc21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6f91c",
    x"020900000000000002aa00000000000000fb337fc31c",
    x"030b00000000000002aafffffffffffff50003e5451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45e01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd328e1c",
    x"070a00000000000002aafffffffffffff8ef3601e81c",
    x"080200000000000002aafffffffffffff6f669e8c61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcbe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6fa1c",
    x"020900000000000002aa00000000000000fb337fbe1c",
    x"030b00000000000002aafffffffffffff50003e5461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf0e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45dc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32881c",
    x"070a00000000000002aafffffffffffff8ef3601e41c",
    x"080200000000000002aafffffffffffff6f669e8c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcb91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6fb1c",
    x"020900000000000002aa00000000000000fb337fb81c",
    x"030b00000000000002aafffffffffffff50003e5471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf0c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32821c",
    x"070a00000000000002aafffffffffffff8ef3601e11c",
    x"080200000000000002aafffffffffffff6f669e8c11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcb51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6fd1c",
    x"020900000000000002aa00000000000000fb337fb31c",
    x"030b00000000000002aafffffffffffff50003e5481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45d51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd327c1c",
    x"070a00000000000002aafffffffffffff8ef3601dd1c",
    x"080200000000000002aafffffffffffff6f669e8bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcb11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6fe1c",
    x"020900000000000002aa00000000000000fb337fad1c",
    x"030b00000000000002aafffffffffffff50003e5491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32761c",
    x"070a00000000000002aafffffffffffff8ef3601da1c",
    x"080200000000000002aafffffffffffff6f669e8bc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dcad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe6ff1c",
    x"020900000000000002aa00000000000000fb337fa71c",
    x"030b00000000000002aafffffffffffff50003e54a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32701c",
    x"070a00000000000002aafffffffffffff8ef3601d61c",
    x"080200000000000002aafffffffffffff6f669e8ba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dca91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7001c",
    x"020900000000000002aa00000000000000fb337fa21c",
    x"030b00000000000002aafffffffffffff50003e54b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45ca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32691c",
    x"070a00000000000002aafffffffffffff8ef3601d21c",
    x"080200000000000002aafffffffffffff6f669e8b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dca41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7011c",
    x"020900000000000002aa00000000000000fb337f9c1c",
    x"030b00000000000002aafffffffffffff50003e54c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcf001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45c61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32631c",
    x"070a00000000000002aafffffffffffff8ef3601cf1c",
    x"080200000000000002aafffffffffffff6f669e8b51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dca01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7021c",
    x"020900000000000002aa00000000000000fb337f971c",
    x"030b00000000000002aafffffffffffff50003e54d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcefe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd325d1c",
    x"070a00000000000002aafffffffffffff8ef3601cb1c",
    x"080200000000000002aafffffffffffff6f669e8b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7031c",
    x"020900000000000002aa00000000000000fb337f911c",
    x"030b00000000000002aafffffffffffff50003e54e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcefb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd32571c",
    x"070a00000000000002aafffffffffffff8ef3601c81c",
    x"080200000000000002aafffffffffffff6f669e8b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266dc981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe7041c",
    x"0209000000000000025a00000000000000fb337f8b1c",
    x"030b000000000000025afffffffffffff50003e54f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dcef91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f45bb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd32511c",
    x"070a000000000000025afffffffffffff8ef3601c41c",
    x"0802000000000000025afffffffffffff6f669e8ae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7051c",
    x"0209000000000000015500000000000000fb337f861c",
    x"030b0000000000000155fffffffffffff50003e5501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcef61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd324b1c",
    x"070a0000000000000155fffffffffffff8ef3601c01c",
    x"08020000000000000155fffffffffffff6f669e8ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dc8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7061c",
    x"0209000000000000031f00000000000000fb337f801c",
    x"030b000000000000031ffffffffffffff50003e5511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcef41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f45b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd32451c",
    x"070a000000000000031ffffffffffffff8ef3601bd1c",
    x"0802000000000000031ffffffffffffff6f669e8a91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dc8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7081c",
    x"020900000000000000ae00000000000000fb337f7b1c",
    x"030b00000000000000aefffffffffffff50003e5521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcef21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f45b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd323e1c",
    x"070a00000000000000aefffffffffffff8ef3601b91c",
    x"080200000000000000aefffffffffffff6f669e8a71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dc871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7091c",
    x"020900000000000001a400000000000000fb337f751c",
    x"030b00000000000001a4fffffffffffff50003e5531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dceef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f45ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd32381c",
    x"070a00000000000001a4fffffffffffff8ef3601b61c",
    x"080200000000000001a4fffffffffffff6f669e8a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266dc831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe70a1c",
    x"0209000000000000019a00000000000000fb337f6f1c",
    x"030b000000000000019afffffffffffff50003e5541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dceed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f45a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd32321c",
    x"070a000000000000019afffffffffffff8ef3601b21c",
    x"0802000000000000019afffffffffffff6f669e8a21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe70b1c",
    x"0209000000000000015500000000000000fb337f6a1c",
    x"030b0000000000000155fffffffffffff50003e5551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dceea1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd322c1c",
    x"070a0000000000000155fffffffffffff8ef3601af1c",
    x"08020000000000000155fffffffffffff6f669e8a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc7a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe70c1c",
    x"0209000000000000015500000000000000fb337f641c",
    x"030b0000000000000155fffffffffffff50003e5561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcee81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32261c",
    x"070a0000000000000155fffffffffffff8ef3601ab1c",
    x"08020000000000000155fffffffffffff6f669e89e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe70d1c",
    x"0209000000000000015500000000000000fb337f5f1c",
    x"030b0000000000000155fffffffffffff50003e5571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcee61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f459d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32201c",
    x"070a0000000000000155fffffffffffff8ef3601a71c",
    x"08020000000000000155fffffffffffff6f669e89b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe70e1c",
    x"0209000000000000015500000000000000fb337f591c",
    x"030b0000000000000155fffffffffffff50003e5581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcee31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f459a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd321a1c",
    x"070a0000000000000155fffffffffffff8ef3601a41c",
    x"08020000000000000155fffffffffffff6f669e8991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe70f1c",
    x"0209000000000000015500000000000000fb337f531c",
    x"030b0000000000000155fffffffffffff50003e5591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcee11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32131c",
    x"070a0000000000000155fffffffffffff8ef3601a01c",
    x"08020000000000000155fffffffffffff6f669e8961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7101c",
    x"0209000000000000015500000000000000fb337f4e1c",
    x"030b0000000000000155fffffffffffff50003e55a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcedf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd320d1c",
    x"070a0000000000000155fffffffffffff8ef36019d1c",
    x"08020000000000000155fffffffffffff6f669e8941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7111c",
    x"0209000000000000015500000000000000fb337f481c",
    x"030b0000000000000155fffffffffffff50003e55b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcedc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f458e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32071c",
    x"070a0000000000000155fffffffffffff8ef3601991c",
    x"08020000000000000155fffffffffffff6f669e8921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7121c",
    x"0209000000000000015500000000000000fb337f431c",
    x"030b0000000000000155fffffffffffff50003e55c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dceda1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f458b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd32011c",
    x"070a0000000000000155fffffffffffff8ef3601951c",
    x"08020000000000000155fffffffffffff6f669e88f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7141c",
    x"0209000000000000015500000000000000fb337f3d1c",
    x"030b0000000000000155fffffffffffff50003e55d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dced71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31fb1c",
    x"070a0000000000000155fffffffffffff8ef3601921c",
    x"08020000000000000155fffffffffffff6f669e88d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7151c",
    x"0209000000000000015500000000000000fb337f371c",
    x"030b0000000000000155fffffffffffff50003e55e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dced51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45831c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31f51c",
    x"070a0000000000000155fffffffffffff8ef36018e1c",
    x"08020000000000000155fffffffffffff6f669e88b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7161c",
    x"0209000000000000015500000000000000fb337f321c",
    x"030b0000000000000155fffffffffffff50003e55f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dced31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31ef1c",
    x"070a0000000000000155fffffffffffff8ef36018b1c",
    x"08020000000000000155fffffffffffff6f669e8881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7171c",
    x"0209000000000000015500000000000000fb337f2c1c",
    x"030b0000000000000155fffffffffffff50003e5601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dced01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f457c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31e91c",
    x"070a0000000000000155fffffffffffff8ef3601871c",
    x"08020000000000000155fffffffffffff6f669e8861c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7181c",
    x"0209000000000000015500000000000000fb337f271c",
    x"030b0000000000000155fffffffffffff50003e5611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcece1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31e21c",
    x"070a0000000000000155fffffffffffff8ef3601841c",
    x"08020000000000000155fffffffffffff6f669e8831c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7191c",
    x"0209000000000000015500000000000000fb337f211c",
    x"030b0000000000000155fffffffffffff50003e5621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcecc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31dc1c",
    x"070a0000000000000155fffffffffffff8ef3601801c",
    x"08020000000000000155fffffffffffff6f669e8811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe71a1c",
    x"0209000000000000015500000000000000fb337f1b1c",
    x"030b0000000000000155fffffffffffff50003e5631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcec91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31d61c",
    x"070a0000000000000155fffffffffffff8ef36017c1c",
    x"08020000000000000155fffffffffffff6f669e87f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe71b1c",
    x"0209000000000000015500000000000000fb337f161c",
    x"030b0000000000000155fffffffffffff50003e5641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcec71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f456d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31d01c",
    x"070a0000000000000155fffffffffffff8ef3601791c",
    x"08020000000000000155fffffffffffff6f669e87c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dc3b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe71c1c",
    x"0209000000000000031f00000000000000fb337f101c",
    x"030b000000000000031ffffffffffffff50003e5651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcec41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f45691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd31ca1c",
    x"070a000000000000031ffffffffffffff8ef3601751c",
    x"0802000000000000031ffffffffffffff6f669e87a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dc371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe71d1c",
    x"020900000000000000ae00000000000000fb337f0b1c",
    x"030b00000000000000aefffffffffffff50003e5661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcec21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f45661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd31c41c",
    x"070a00000000000000aefffffffffffff8ef3601721c",
    x"080200000000000000aefffffffffffff6f669e8771c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dc331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe71f1c",
    x"020900000000000001a400000000000000fb337f051c",
    x"030b00000000000001a4fffffffffffff50003e5671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcec01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f45621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd31be1c",
    x"070a00000000000001a4fffffffffffff8ef36016e1c",
    x"080200000000000001a4fffffffffffff6f669e8751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266dc2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe7201c",
    x"0209000000000000015600000000000000fb337f001c",
    x"030b0000000000000156fffffffffffff50003e5681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dcebd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f455e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd31b71c",
    x"070a0000000000000156fffffffffffff8ef36016a1c",
    x"08020000000000000156fffffffffffff6f669e8731c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dc2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7211c",
    x"0209000000000000015500000000000000fb337efa1c",
    x"030b0000000000000155fffffffffffff50003e5691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcebb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f455b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31b11c",
    x"070a0000000000000155fffffffffffff8ef3601671c",
    x"08020000000000000155fffffffffffff6f669e8701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266dc261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe7221c",
    x"0209000000000000029a00000000000000fb337ef41c",
    x"030b000000000000029afffffffffffff50003e56a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dceb81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f45571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd31ab1c",
    x"070a000000000000029afffffffffffff8ef3601631c",
    x"0802000000000000029afffffffffffff6f669e86e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7231c",
    x"020900000000000002aa00000000000000fb337eef1c",
    x"030b00000000000002aafffffffffffff50003e56b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dceb61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31a51c",
    x"070a00000000000002aafffffffffffff8ef3601601c",
    x"080200000000000002aafffffffffffff6f669e86c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7241c",
    x"020900000000000002aa00000000000000fb337ee91c",
    x"030b00000000000002aafffffffffffff50003e56c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dceb41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f454f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd319f1c",
    x"070a00000000000002aafffffffffffff8ef36015c1c",
    x"080200000000000002aafffffffffffff6f669e8691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7251c",
    x"020900000000000002aa00000000000000fb337ee41c",
    x"030b00000000000002aafffffffffffff50003e56d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dceb11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f454c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31991c",
    x"070a00000000000002aafffffffffffff8ef3601591c",
    x"080200000000000002aafffffffffffff6f669e8671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7261c",
    x"020900000000000002aa00000000000000fb337ede1c",
    x"030b00000000000002aafffffffffffff50003e56e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dceaf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31931c",
    x"070a00000000000002aafffffffffffff8ef3601551c",
    x"080200000000000002aafffffffffffff6f669e8641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7271c",
    x"020900000000000002aa00000000000000fb337ed81c",
    x"030b00000000000002aafffffffffffff50003e56f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcead1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd318c1c",
    x"070a00000000000002aafffffffffffff8ef3601511c",
    x"080200000000000002aafffffffffffff6f669e8621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc0d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7281c",
    x"020900000000000002aa00000000000000fb337ed31c",
    x"030b00000000000002aafffffffffffff50003e5701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dceaa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31861c",
    x"070a00000000000002aafffffffffffff8ef36014e1c",
    x"080200000000000002aafffffffffffff6f669e8601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe72a1c",
    x"020900000000000002aa00000000000000fb337ecd1c",
    x"030b00000000000002aafffffffffffff50003e5711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcea81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f453d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31801c",
    x"070a00000000000002aafffffffffffff8ef36014a1c",
    x"080200000000000002aafffffffffffff6f669e85d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe72b1c",
    x"020900000000000002aa00000000000000fb337ec81c",
    x"030b00000000000002aafffffffffffff50003e5721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcea51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd317a1c",
    x"070a00000000000002aafffffffffffff8ef3601471c",
    x"080200000000000002aafffffffffffff6f669e85b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dc011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe72c1c",
    x"020900000000000002aa00000000000000fb337ec21c",
    x"030b00000000000002aafffffffffffff50003e5731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcea31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31741c",
    x"070a00000000000002aafffffffffffff8ef3601431c",
    x"080200000000000002aafffffffffffff6f669e8591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbfc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe72d1c",
    x"020900000000000002aa00000000000000fb337ebc1c",
    x"030b00000000000002aafffffffffffff50003e5741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcea11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd316e1c",
    x"070a00000000000002aafffffffffffff8ef36013f1c",
    x"080200000000000002aafffffffffffff6f669e8561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbf81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe72e1c",
    x"020900000000000002aa00000000000000fb337eb71c",
    x"030b00000000000002aafffffffffffff50003e5751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce9e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f452e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31681c",
    x"070a00000000000002aafffffffffffff8ef36013c1c",
    x"080200000000000002aafffffffffffff6f669e8541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbf41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe72f1c",
    x"020900000000000002aa00000000000000fb337eb11c",
    x"030b00000000000002aafffffffffffff50003e5771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce9c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f452a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31611c",
    x"070a00000000000002aafffffffffffff8ef3601381c",
    x"080200000000000002aafffffffffffff6f669e8511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266dbf01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe7301c",
    x"0209000000000000026a00000000000000fb337eac1c",
    x"030b000000000000026afffffffffffff50003e5781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dce991c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f45271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026affffffffffffff04cd315b1c",
    x"070a000000000000026afffffffffffff8ef3601351c",
    x"0802000000000000026afffffffffffff6f669e84f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dbec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7311c",
    x"0209000000000000015500000000000000fb337ea61c",
    x"030b0000000000000155fffffffffffff50003e5791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f45231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd31551c",
    x"070a0000000000000155fffffffffffff8ef3601311c",
    x"08020000000000000155fffffffffffff6f669e84d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266dbe71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7321c",
    x"0209000000000000031f00000000000000fb337ea01c",
    x"030b000000000000031ffffffffffffff50003e57a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dce951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f451f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd314f1c",
    x"070a000000000000031ffffffffffffff8ef36012d1c",
    x"0802000000000000031ffffffffffffff6f669e84a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dbe31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7331c",
    x"020900000000000000ae00000000000000fb337e9b1c",
    x"030b00000000000000aefffffffffffff50003e57b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dce921c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f451c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd31491c",
    x"070a00000000000000aefffffffffffff8ef36012a1c",
    x"080200000000000000aefffffffffffff6f669e8481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dbdf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7341c",
    x"020900000000000001a400000000000000fb337e951c",
    x"030b00000000000001a4fffffffffffff50003e57c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dce901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f45181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd31431c",
    x"070a00000000000001a4fffffffffffff8ef3601261c",
    x"080200000000000001a4fffffffffffff6f669e8461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266dbdb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe7361c",
    x"0209000000000000025600000000000000fb337e901c",
    x"030b0000000000000256fffffffffffff50003e57d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dce8e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f45141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd313d1c",
    x"070a0000000000000256fffffffffffff8ef3601231c",
    x"08020000000000000256fffffffffffff6f669e8431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbd71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7371c",
    x"020900000000000002aa00000000000000fb337e8a1c",
    x"030b00000000000002aafffffffffffff50003e57e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce8b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45101c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31361c",
    x"070a00000000000002aafffffffffffff8ef36011f1c",
    x"080200000000000002aafffffffffffff6f669e8411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbd21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7381c",
    x"020900000000000002aa00000000000000fb337e841c",
    x"030b00000000000002aafffffffffffff50003e57f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f450d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31301c",
    x"070a00000000000002aafffffffffffff8ef36011c1c",
    x"080200000000000002aafffffffffffff6f669e83e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7391c",
    x"020900000000000002aa00000000000000fb337e7f1c",
    x"030b00000000000002aafffffffffffff50003e5801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd312a1c",
    x"070a00000000000002aafffffffffffff8ef3601181c",
    x"080200000000000002aafffffffffffff6f669e83c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe73a1c",
    x"020900000000000002aa00000000000000fb337e791c",
    x"030b00000000000002aafffffffffffff50003e5811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31241c",
    x"070a00000000000002aafffffffffffff8ef3601141c",
    x"080200000000000002aafffffffffffff6f669e83a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbc61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe73b1c",
    x"020900000000000002aa00000000000000fb337e741c",
    x"030b00000000000002aafffffffffffff50003e5821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f45021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd311e1c",
    x"070a00000000000002aafffffffffffff8ef3601111c",
    x"080200000000000002aafffffffffffff6f669e8371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbc21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe73c1c",
    x"020900000000000002aa00000000000000fb337e6e1c",
    x"030b00000000000002aafffffffffffff50003e5831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce7f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44fe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31181c",
    x"070a00000000000002aafffffffffffff8ef36010d1c",
    x"080200000000000002aafffffffffffff6f669e8351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbbe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe73d1c",
    x"020900000000000002aa00000000000000fb337e691c",
    x"030b00000000000002aafffffffffffff50003e5841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce7d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44fa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31121c",
    x"070a00000000000002aafffffffffffff8ef36010a1c",
    x"080200000000000002aafffffffffffff6f669e8321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbb91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe73e1c",
    x"020900000000000002aa00000000000000fb337e631c",
    x"030b00000000000002aafffffffffffff50003e5851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce7a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44f61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd310b1c",
    x"070a00000000000002aafffffffffffff8ef3601061c",
    x"080200000000000002aafffffffffffff6f669e8301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbb51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe73f1c",
    x"020900000000000002aa00000000000000fb337e5d1c",
    x"030b00000000000002aafffffffffffff50003e5861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44f31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd31051c",
    x"070a00000000000002aafffffffffffff8ef3601021c",
    x"080200000000000002aafffffffffffff6f669e82e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbb11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7411c",
    x"020900000000000002aa00000000000000fb337e581c",
    x"030b00000000000002aafffffffffffff50003e5871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44ef1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30ff1c",
    x"070a00000000000002aafffffffffffff8ef3600ff1c",
    x"080200000000000002aafffffffffffff6f669e82b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dbad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7421c",
    x"020900000000000002aa00000000000000fb337e521c",
    x"030b00000000000002aafffffffffffff50003e5881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30f91c",
    x"070a00000000000002aafffffffffffff8ef3600fb1c",
    x"080200000000000002aafffffffffffff6f669e8291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dba91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7431c",
    x"020900000000000002aa00000000000000fb337e4d1c",
    x"030b00000000000002aafffffffffffff50003e5891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44e81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30f31c",
    x"070a00000000000002aafffffffffffff8ef3600f81c",
    x"080200000000000002aafffffffffffff6f669e8271c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dba41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7441c",
    x"020900000000000002aa00000000000000fb337e471c",
    x"030b00000000000002aafffffffffffff50003e58a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce6f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44e41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30ed1c",
    x"070a00000000000002aafffffffffffff8ef3600f41c",
    x"080200000000000002aafffffffffffff6f669e8241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266dba01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7451c",
    x"020900000000000002aa00000000000000fb337e411c",
    x"030b00000000000002aafffffffffffff50003e58b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce6c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44e01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30e71c",
    x"070a00000000000002aafffffffffffff8ef3600f01c",
    x"080200000000000002aafffffffffffff6f669e8221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266db9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe7461c",
    x"0209000000000000029a00000000000000fb337e3c1c",
    x"030b000000000000029afffffffffffff50003e58c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dce6a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f44dd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd30e01c",
    x"070a000000000000029afffffffffffff8ef3600ed1c",
    x"0802000000000000029afffffffffffff6f669e81f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7471c",
    x"020900000000000002aa00000000000000fb337e361c",
    x"030b00000000000002aafffffffffffff50003e58d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30da1c",
    x"070a00000000000002aafffffffffffff8ef3600e91c",
    x"080200000000000002aafffffffffffff6f669e81d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266db941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7481c",
    x"0209000000000000031f00000000000000fb337e311c",
    x"030b000000000000031ffffffffffffff50003e58e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dce651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f44d51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd30d41c",
    x"070a000000000000031ffffffffffffff8ef3600e61c",
    x"0802000000000000031ffffffffffffff6f669e81b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266db8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7491c",
    x"020900000000000000ae00000000000000fb337e2b1c",
    x"030b00000000000000aefffffffffffff50003e58f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dce631c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f44d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd30ce1c",
    x"070a00000000000000aefffffffffffff8ef3600e21c",
    x"080200000000000000aefffffffffffff6f669e8181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266db8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe74a1c",
    x"020900000000000001a400000000000000fb337e251c",
    x"030b00000000000001a4fffffffffffff50003e5901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dce601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f44ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd30c81c",
    x"070a00000000000001a4fffffffffffff8ef3600de1c",
    x"080200000000000001a4fffffffffffff6f669e8161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266db871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe74c1c",
    x"0209000000000000029600000000000000fb337e201c",
    x"030b0000000000000296fffffffffffff50003e5911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dce5e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f44ca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd30c21c",
    x"070a0000000000000296fffffffffffff8ef3600db1c",
    x"08020000000000000296fffffffffffff6f669e8141c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe74d1c",
    x"020900000000000002aa00000000000000fb337e1a1c",
    x"030b00000000000002aafffffffffffff50003e5921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce5b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44c61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30bc1c",
    x"070a00000000000002aafffffffffffff8ef3600d71c",
    x"080200000000000002aafffffffffffff6f669e8111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266db7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe74e1c",
    x"020900000000000002a900000000000000fb337e151c",
    x"030b00000000000002a9fffffffffffff50003e5931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a9fffffffffffff4099dce591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f44c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd30b51c",
    x"070a00000000000002a9fffffffffffff8ef3600d41c",
    x"080200000000000002a9fffffffffffff6f669e80f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db7a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe74f1c",
    x"020900000000000002aa00000000000000fb337e0f1c",
    x"030b00000000000002aafffffffffffff50003e5941c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30af1c",
    x"070a00000000000002aafffffffffffff8ef3600d01c",
    x"080200000000000002aafffffffffffff6f669e80c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7501c",
    x"020900000000000002aa00000000000000fb337e091c",
    x"030b00000000000002aafffffffffffff50003e5951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44bb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30a91c",
    x"070a00000000000002aafffffffffffff8ef3600cd1c",
    x"080200000000000002aafffffffffffff6f669e80a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7511c",
    x"020900000000000002aa00000000000000fb337e041c",
    x"030b00000000000002aafffffffffffff50003e5961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44b81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30a31c",
    x"070a00000000000002aafffffffffffff8ef3600c91c",
    x"080200000000000002aafffffffffffff6f669e8081c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7521c",
    x"020900000000000002aa00000000000000fb337dfe1c",
    x"030b00000000000002aafffffffffffff50003e5971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce4f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd309d1c",
    x"070a00000000000002aafffffffffffff8ef3600c51c",
    x"080200000000000002aafffffffffffff6f669e8051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7531c",
    x"020900000000000002aa00000000000000fb337df91c",
    x"030b00000000000002aafffffffffffff50003e5981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce4d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30971c",
    x"070a00000000000002aafffffffffffff8ef3600c21c",
    x"080200000000000002aafffffffffffff6f669e8031c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7541c",
    x"020900000000000002aa00000000000000fb337df31c",
    x"030b00000000000002aafffffffffffff50003e5991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce4b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30911c",
    x"070a00000000000002aafffffffffffff8ef3600be1c",
    x"080200000000000002aafffffffffffff6f669e8001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7551c",
    x"020900000000000002aa00000000000000fb337ded1c",
    x"030b00000000000002aafffffffffffff50003e59a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44a91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd308a1c",
    x"070a00000000000002aafffffffffffff8ef3600bb1c",
    x"080200000000000002aafffffffffffff6f669e7fe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7571c",
    x"020900000000000002aa00000000000000fb337de81c",
    x"030b00000000000002aafffffffffffff50003e59b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30841c",
    x"070a00000000000002aafffffffffffff8ef3600b71c",
    x"080200000000000002aafffffffffffff6f669e7fc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7581c",
    x"020900000000000002aa00000000000000fb337de21c",
    x"030b00000000000002aafffffffffffff50003e59c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd307e1c",
    x"070a00000000000002aafffffffffffff8ef3600b31c",
    x"080200000000000002aafffffffffffff6f669e7f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7591c",
    x"020900000000000002aa00000000000000fb337ddd1c",
    x"030b00000000000002aafffffffffffff50003e59d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f449e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30781c",
    x"070a00000000000002aafffffffffffff8ef3600b01c",
    x"080200000000000002aafffffffffffff6f669e7f71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe75a1c",
    x"020900000000000002aa00000000000000fb337dd71c",
    x"030b00000000000002aafffffffffffff50003e59e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce3f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f449a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd30721c",
    x"070a00000000000002aafffffffffffff8ef3600ac1c",
    x"080200000000000002aafffffffffffff6f669e7f51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266db4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe75b1c",
    x"020900000000000002aa00000000000000fb337dd11c",
    x"030b00000000000002aafffffffffffff50003e59f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce3c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd306c1c",
    x"070a00000000000002aafffffffffffff8ef3600a91c",
    x"080200000000000002aafffffffffffff6f669e7f21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266db481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe75c1c",
    x"0209000000000000015a00000000000000fb337dcc1c",
    x"030b000000000000015afffffffffffff50003e5a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dce3a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f44921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd30661c",
    x"070a000000000000015afffffffffffff8ef3600a51c",
    x"0802000000000000015afffffffffffff6f669e7f01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe75d1c",
    x"0209000000000000015500000000000000fb337dc61c",
    x"030b0000000000000155fffffffffffff50003e5a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f448f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd305f1c",
    x"070a0000000000000155fffffffffffff8ef3600a11c",
    x"08020000000000000155fffffffffffff6f669e7ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266db401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe75e1c",
    x"0209000000000000031f00000000000000fb337dc11c",
    x"030b000000000000031ffffffffffffff50003e5a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dce351c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f448b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd30591c",
    x"070a000000000000031ffffffffffffff8ef36009e1c",
    x"0802000000000000031ffffffffffffff6f669e7eb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266db3b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe75f1c",
    x"020900000000000000ae00000000000000fb337dbb1c",
    x"030b00000000000000aefffffffffffff50003e5a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dce331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f44871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd30531c",
    x"070a00000000000000aefffffffffffff8ef36009a1c",
    x"080200000000000000aefffffffffffff6f669e7e91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266db371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7601c",
    x"020900000000000001a400000000000000fb337db51c",
    x"030b00000000000001a4fffffffffffff50003e5a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dce301c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f44841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd304d1c",
    x"070a00000000000001a4fffffffffffff8ef3600971c",
    x"080200000000000001a4fffffffffffff6f669e7e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266db331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe7621c",
    x"0209000000000000019600000000000000fb337db01c",
    x"030b0000000000000196fffffffffffff50003e5a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dce2e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f44801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000196ffffffffffffff04cd30471c",
    x"070a0000000000000196fffffffffffff8ef3600931c",
    x"08020000000000000196fffffffffffff6f669e7e41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7631c",
    x"0209000000000000015500000000000000fb337daa1c",
    x"030b0000000000000155fffffffffffff50003e5a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce2c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f447c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30411c",
    x"070a0000000000000155fffffffffffff8ef36008f1c",
    x"08020000000000000155fffffffffffff6f669e7e21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7641c",
    x"0209000000000000015500000000000000fb337da51c",
    x"030b0000000000000155fffffffffffff50003e5a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce291c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd303b1c",
    x"070a0000000000000155fffffffffffff8ef36008c1c",
    x"08020000000000000155fffffffffffff6f669e7df1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7651c",
    x"0209000000000000015500000000000000fb337d9f1c",
    x"030b0000000000000155fffffffffffff50003e5a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30351c",
    x"070a0000000000000155fffffffffffff8ef3600881c",
    x"08020000000000000155fffffffffffff6f669e7dd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7661c",
    x"0209000000000000015500000000000000fb337d9a1c",
    x"030b0000000000000155fffffffffffff50003e5a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd302e1c",
    x"070a0000000000000155fffffffffffff8ef3600851c",
    x"08020000000000000155fffffffffffff6f669e7da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7671c",
    x"0209000000000000015500000000000000fb337d941c",
    x"030b0000000000000155fffffffffffff50003e5aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f446d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30281c",
    x"070a0000000000000155fffffffffffff8ef3600811c",
    x"08020000000000000155fffffffffffff6f669e7d81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7681c",
    x"0209000000000000015500000000000000fb337d8e1c",
    x"030b0000000000000155fffffffffffff50003e5ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f446a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30221c",
    x"070a0000000000000155fffffffffffff8ef36007d1c",
    x"08020000000000000155fffffffffffff6f669e7d61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7691c",
    x"0209000000000000015500000000000000fb337d891c",
    x"030b0000000000000155fffffffffffff50003e5ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce1d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd301c1c",
    x"070a0000000000000155fffffffffffff8ef36007a1c",
    x"08020000000000000155fffffffffffff6f669e7d31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe76a1c",
    x"0209000000000000015500000000000000fb337d831c",
    x"030b0000000000000155fffffffffffff50003e5ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce1b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30161c",
    x"070a0000000000000155fffffffffffff8ef3600761c",
    x"08020000000000000155fffffffffffff6f669e7d11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db0d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe76b1c",
    x"0209000000000000015500000000000000fb337d7e1c",
    x"030b0000000000000155fffffffffffff50003e5ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f445f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30101c",
    x"070a0000000000000155fffffffffffff8ef3600731c",
    x"08020000000000000155fffffffffffff6f669e7ce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe76d1c",
    x"0209000000000000015500000000000000fb337d781c",
    x"030b0000000000000155fffffffffffff50003e5af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f445b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd300a1c",
    x"070a0000000000000155fffffffffffff8ef36006f1c",
    x"08020000000000000155fffffffffffff6f669e7cc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe76e1c",
    x"0209000000000000015500000000000000fb337d721c",
    x"030b0000000000000155fffffffffffff50003e5b01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd30031c",
    x"070a0000000000000155fffffffffffff8ef36006c1c",
    x"08020000000000000155fffffffffffff6f669e7ca1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266db011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe76f1c",
    x"0209000000000000015500000000000000fb337d6d1c",
    x"030b0000000000000155fffffffffffff50003e5b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ffd1c",
    x"070a0000000000000155fffffffffffff8ef3600681c",
    x"08020000000000000155fffffffffffff6f669e7c71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dafd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7701c",
    x"0209000000000000015500000000000000fb337d671c",
    x"030b0000000000000155fffffffffffff50003e5b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce0f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ff71c",
    x"070a0000000000000155fffffffffffff8ef3600641c",
    x"08020000000000000155fffffffffffff6f669e7c51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266daf81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7711c",
    x"0209000000000000015500000000000000fb337d621c",
    x"030b0000000000000155fffffffffffff50003e5b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dce0d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f444c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ff11c",
    x"070a0000000000000155fffffffffffff8ef3600611c",
    x"08020000000000000155fffffffffffff6f669e7c31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266daf41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbe7721c",
    x"020900000000000002a500000000000000fb337d5c1c",
    x"030b00000000000002a5fffffffffffff50003e5b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dce0a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f44481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd2feb1c",
    x"070a00000000000002a5fffffffffffff8ef36005d1c",
    x"080200000000000002a5fffffffffffff6f669e7c01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266daf01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7731c",
    x"020900000000000002aa00000000000000fb337d561c",
    x"030b00000000000002aafffffffffffff50003e5b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dce081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f44451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2fe51c",
    x"070a00000000000002aafffffffffffff8ef36005a1c",
    x"080200000000000002aafffffffffffff6f669e7be1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266daec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7741c",
    x"0209000000000000031f00000000000000fb337d511c",
    x"030b000000000000031ffffffffffffff50003e5b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dce051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f44411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2fdf1c",
    x"070a000000000000031ffffffffffffff8ef3600561c",
    x"0802000000000000031ffffffffffffff6f669e7bb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266dae81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7751c",
    x"020900000000000000ae00000000000000fb337d4b1c",
    x"030b00000000000000aefffffffffffff50003e5b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dce031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f443d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2fd81c",
    x"070a00000000000000aefffffffffffff8ef3600521c",
    x"080200000000000000aefffffffffffff6f669e7b91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266dae31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7761c",
    x"020900000000000001a400000000000000fb337d461c",
    x"030b00000000000001a4fffffffffffff50003e5b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dce011c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f443a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2fd21c",
    x"070a00000000000001a4fffffffffffff8ef36004f1c",
    x"080200000000000001a4fffffffffffff6f669e7b71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266dadf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbe7771c",
    x"020900000000000002a600000000000000fb337d401c",
    x"030b00000000000002a6fffffffffffff50003e5b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dcdfe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f44361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd2fcc1c",
    x"070a00000000000002a6fffffffffffff8ef36004b1c",
    x"080200000000000002a6fffffffffffff6f669e7b41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266dadb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe7791c",
    x"0209000000000000016a00000000000000fb337d3a1c",
    x"030b000000000000016afffffffffffff50003e5ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcdfc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f44321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd2fc61c",
    x"070a000000000000016afffffffffffff8ef3600481c",
    x"0802000000000000016afffffffffffff6f669e7b21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266dad71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe77a1c",
    x"0209000000000000016900000000000000fb337d351c",
    x"030b0000000000000169fffffffffffff50003e5bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dcdf91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001690000000000000b072f442f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd2fc01c",
    x"070a0000000000000169fffffffffffff8ef3600441c",
    x"08020000000000000169fffffffffffff6f669e7af1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dad31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe77b1c",
    x"0209000000000000015500000000000000fb337d2f1c",
    x"030b0000000000000155fffffffffffff50003e5bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdf71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f442b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2fba1c",
    x"070a0000000000000155fffffffffffff8ef3600401c",
    x"08020000000000000155fffffffffffff6f669e7ad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dace1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe77c1c",
    x"0209000000000000015500000000000000fb337d2a1c",
    x"030b0000000000000155fffffffffffff50003e5bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdf51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2fb41c",
    x"070a0000000000000155fffffffffffff8ef36003d1c",
    x"08020000000000000155fffffffffffff6f669e7ab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266daca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe77d1c",
    x"0209000000000000015500000000000000fb337d241c",
    x"030b0000000000000155fffffffffffff50003e5be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdf21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2fad1c",
    x"070a0000000000000155fffffffffffff8ef3600391c",
    x"08020000000000000155fffffffffffff6f669e7a81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dac61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe77e1c",
    x"0209000000000000015500000000000000fb337d1e1c",
    x"030b0000000000000155fffffffffffff50003e5bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdf01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2fa71c",
    x"070a0000000000000155fffffffffffff8ef3600361c",
    x"08020000000000000155fffffffffffff6f669e7a61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dac21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe77f1c",
    x"0209000000000000015500000000000000fb337d191c",
    x"030b0000000000000155fffffffffffff50003e5c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcded1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f441c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2fa11c",
    x"070a0000000000000155fffffffffffff8ef3600321c",
    x"08020000000000000155fffffffffffff6f669e7a41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dabe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7801c",
    x"0209000000000000015500000000000000fb337d131c",
    x"030b0000000000000155fffffffffffff50003e5c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdeb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f9b1c",
    x"070a0000000000000155fffffffffffff8ef36002e1c",
    x"08020000000000000155fffffffffffff6f669e7a11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dab91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7811c",
    x"0209000000000000015500000000000000fb337d0e1c",
    x"030b0000000000000155fffffffffffff50003e5c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcde91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f951c",
    x"070a0000000000000155fffffffffffff8ef36002b1c",
    x"08020000000000000155fffffffffffff6f669e79f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dab51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7821c",
    x"0209000000000000015500000000000000fb337d081c",
    x"030b0000000000000155fffffffffffff50003e5c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcde61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f8f1c",
    x"070a0000000000000155fffffffffffff8ef3600271c",
    x"08020000000000000155fffffffffffff6f669e79c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266dab11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7841c",
    x"0209000000000000015500000000000000fb337d021c",
    x"030b0000000000000155fffffffffffff50003e5c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcde41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f440d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f891c",
    x"070a0000000000000155fffffffffffff8ef3600241c",
    x"08020000000000000155fffffffffffff6f669e79a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266daad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7851c",
    x"0209000000000000015500000000000000fb337cfd1c",
    x"030b0000000000000155fffffffffffff50003e5c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcde21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f440a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f821c",
    x"070a0000000000000155fffffffffffff8ef3600201c",
    x"08020000000000000155fffffffffffff6f669e7981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266daa91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7861c",
    x"0209000000000000015500000000000000fb337cf71c",
    x"030b0000000000000155fffffffffffff50003e5c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcddf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f7c1c",
    x"070a0000000000000155fffffffffffff8ef36001c1c",
    x"08020000000000000155fffffffffffff6f669e7951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266daa41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7871c",
    x"0209000000000000015500000000000000fb337cf21c",
    x"030b0000000000000155fffffffffffff50003e5c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcddd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f44021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f761c",
    x"070a0000000000000155fffffffffffff8ef3600191c",
    x"08020000000000000155fffffffffffff6f669e7931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266daa01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7881c",
    x"0209000000000000015500000000000000fb337cec1c",
    x"030b0000000000000155fffffffffffff50003e5c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdda1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43fe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f701c",
    x"070a0000000000000155fffffffffffff8ef3600151c",
    x"08020000000000000155fffffffffffff6f669e7911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7891c",
    x"0209000000000000015500000000000000fb337ce61c",
    x"030b0000000000000155fffffffffffff50003e5c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdd81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f6a1c",
    x"070a0000000000000155fffffffffffff8ef3600121c",
    x"08020000000000000155fffffffffffff6f669e78e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266da981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe78a1c",
    x"0209000000000000031f00000000000000fb337ce11c",
    x"030b000000000000031ffffffffffffff50003e5cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcdd61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f43f71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2f641c",
    x"070a000000000000031ffffffffffffff8ef36000e1c",
    x"0802000000000000031ffffffffffffff6f669e78c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266da941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe78b1c",
    x"020900000000000000ae00000000000000fb337cdb1c",
    x"030b00000000000000aefffffffffffff50003e5cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcdd31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f43f31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2f5e1c",
    x"070a00000000000000aefffffffffffff8ef36000a1c",
    x"080200000000000000aefffffffffffff6f669e7891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266da8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe78c1c",
    x"020900000000000001a400000000000000fb337cd61c",
    x"030b00000000000001a4fffffffffffff50003e5cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcdd11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f43f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2f571c",
    x"070a00000000000001a4fffffffffffff8ef3600071c",
    x"080200000000000001a4fffffffffffff6f669e7871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266da8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe78d1c",
    x"020900000000000001a600000000000000fb337cd01c",
    x"030b00000000000001a6fffffffffffff50003e5ce1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dcdce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f43ec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd2f511c",
    x"070a00000000000001a6fffffffffffff8ef3600031c",
    x"080200000000000001a6fffffffffffff6f669e7851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe78f1c",
    x"0209000000000000015500000000000000fb337cca1c",
    x"030b0000000000000155fffffffffffff50003e5cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdcc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43e81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f4b1c",
    x"070a0000000000000155fffffffffffff8ef3600001c",
    x"08020000000000000155fffffffffffff6f669e7821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7901c",
    x"0209000000000000015500000000000000fb337cc51c",
    x"030b0000000000000155fffffffffffff50003e5d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43e51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f451c",
    x"070a0000000000000155fffffffffffff8ef35fffc1c",
    x"08020000000000000155fffffffffffff6f669e7801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7911c",
    x"0209000000000000015500000000000000fb337cbf1c",
    x"030b0000000000000155fffffffffffff50003e5d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdc71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43e11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f3f1c",
    x"070a0000000000000155fffffffffffff8ef35fff81c",
    x"08020000000000000155fffffffffffff6f669e77d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da7a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7921c",
    x"0209000000000000015500000000000000fb337cba1c",
    x"030b0000000000000155fffffffffffff50003e5d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdc51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43dd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f391c",
    x"070a0000000000000155fffffffffffff8ef35fff51c",
    x"08020000000000000155fffffffffffff6f669e77b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7931c",
    x"0209000000000000015500000000000000fb337cb41c",
    x"030b0000000000000155fffffffffffff50003e5d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdc21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f331c",
    x"070a0000000000000155fffffffffffff8ef35fff11c",
    x"08020000000000000155fffffffffffff6f669e7791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7941c",
    x"0209000000000000015500000000000000fb337caf1c",
    x"030b0000000000000155fffffffffffff50003e5d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdc01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43d61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f2c1c",
    x"070a0000000000000155fffffffffffff8ef35ffee1c",
    x"08020000000000000155fffffffffffff6f669e7761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7951c",
    x"0209000000000000015500000000000000fb337ca91c",
    x"030b0000000000000155fffffffffffff50003e5d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdbe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43d21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f261c",
    x"070a0000000000000155fffffffffffff8ef35ffea1c",
    x"08020000000000000155fffffffffffff6f669e7741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7961c",
    x"0209000000000000015500000000000000fb337ca31c",
    x"030b0000000000000155fffffffffffff50003e5d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdbb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f201c",
    x"070a0000000000000155fffffffffffff8ef35ffe61c",
    x"08020000000000000155fffffffffffff6f669e7721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7971c",
    x"0209000000000000015500000000000000fb337c9e1c",
    x"030b0000000000000155fffffffffffff50003e5d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdb91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43cb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f1a1c",
    x"070a0000000000000155fffffffffffff8ef35ffe31c",
    x"08020000000000000155fffffffffffff6f669e76f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7981c",
    x"0209000000000000015500000000000000fb337c981c",
    x"030b0000000000000155fffffffffffff50003e5d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdb61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43c71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f141c",
    x"070a0000000000000155fffffffffffff8ef35ffdf1c",
    x"08020000000000000155fffffffffffff6f669e76d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe79a1c",
    x"0209000000000000015500000000000000fb337c931c",
    x"030b0000000000000155fffffffffffff50003e5d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdb41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f0e1c",
    x"070a0000000000000155fffffffffffff8ef35ffdc1c",
    x"08020000000000000155fffffffffffff6f669e76a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe79b1c",
    x"0209000000000000015500000000000000fb337c8d1c",
    x"030b0000000000000155fffffffffffff50003e5da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdb21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43c01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f071c",
    x"070a0000000000000155fffffffffffff8ef35ffd81c",
    x"08020000000000000155fffffffffffff6f669e7681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe79c1c",
    x"0209000000000000015500000000000000fb337c871c",
    x"030b0000000000000155fffffffffffff50003e5db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdaf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43bc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2f011c",
    x"070a0000000000000155fffffffffffff8ef35ffd41c",
    x"08020000000000000155fffffffffffff6f669e7661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe79d1c",
    x"0209000000000000015500000000000000fb337c821c",
    x"030b0000000000000155fffffffffffff50003e5dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcdad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43b81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2efb1c",
    x"070a0000000000000155fffffffffffff8ef35ffd11c",
    x"08020000000000000155fffffffffffff6f669e7631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266da4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe79e1c",
    x"0209000000000000029500000000000000fb337c7c1c",
    x"030b0000000000000295fffffffffffff50003e5dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcdaa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f43b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2ef51c",
    x"070a0000000000000295fffffffffffff8ef35ffcd1c",
    x"08020000000000000295fffffffffffff6f669e7611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266da481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe79f1c",
    x"020900000000000002aa00000000000000fb337c771c",
    x"030b00000000000002aafffffffffffff50003e5de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcda81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43b11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2eef1c",
    x"070a00000000000002aafffffffffffff8ef35ffca1c",
    x"080200000000000002aafffffffffffff6f669e75e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266da441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7a01c",
    x"0209000000000000031f00000000000000fb337c711c",
    x"030b000000000000031ffffffffffffff50003e5df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcda61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f43ad1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2ee91c",
    x"070a000000000000031ffffffffffffff8ef35ffc61c",
    x"0802000000000000031ffffffffffffff6f669e75c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266da401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7a11c",
    x"020900000000000000ae00000000000000fb337c6b1c",
    x"030b00000000000000aefffffffffffff50003e5e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcda31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f43a91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2ee31c",
    x"070a00000000000000aefffffffffffff8ef35ffc21c",
    x"080200000000000000aefffffffffffff6f669e75a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266da3c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7a21c",
    x"020900000000000001a400000000000000fb337c661c",
    x"030b00000000000001a4fffffffffffff50003e5e11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcda11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f43a61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2edc1c",
    x"070a00000000000001a4fffffffffffff8ef35ffbf1c",
    x"080200000000000001a4fffffffffffff6f669e7571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266da371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe7a31c",
    x"0209000000000000016600000000000000fb337c601c",
    x"030b0000000000000166fffffffffffff50003e5e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dcd9e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f43a21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd2ed61c",
    x"070a0000000000000166fffffffffffff8ef35ffbb1c",
    x"08020000000000000166fffffffffffff6f669e7551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266da331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe7a51c",
    x"0209000000000000029500000000000000fb337c5b1c",
    x"030b0000000000000295fffffffffffff50003e5e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcd9c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f439e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2ed01c",
    x"070a0000000000000295fffffffffffff8ef35ffb81c",
    x"08020000000000000295fffffffffffff6f669e7531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266da2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe7a61c",
    x"0209000000000000015900000000000000fb337c551c",
    x"030b0000000000000159fffffffffffff50003e5e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcd9a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f439b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd2eca1c",
    x"070a0000000000000159fffffffffffff8ef35ffb41c",
    x"08020000000000000159fffffffffffff6f669e7501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7a71c",
    x"0209000000000000015500000000000000fb337c4f1c",
    x"030b0000000000000155fffffffffffff50003e5e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43971c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ec41c",
    x"070a0000000000000155fffffffffffff8ef35ffb01c",
    x"08020000000000000155fffffffffffff6f669e74e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7a81c",
    x"0209000000000000015500000000000000fb337c4a1c",
    x"030b0000000000000155fffffffffffff50003e5e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ebe1c",
    x"070a0000000000000155fffffffffffff8ef35ffad1c",
    x"08020000000000000155fffffffffffff6f669e74b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7a91c",
    x"0209000000000000015500000000000000fb337c441c",
    x"030b0000000000000155fffffffffffff50003e5e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f438f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2eb81c",
    x"070a0000000000000155fffffffffffff8ef35ffa91c",
    x"08020000000000000155fffffffffffff6f669e7491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7aa1c",
    x"0209000000000000015500000000000000fb337c3f1c",
    x"030b0000000000000155fffffffffffff50003e5e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f438c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2eb11c",
    x"070a0000000000000155fffffffffffff8ef35ffa61c",
    x"08020000000000000155fffffffffffff6f669e7471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7ab1c",
    x"0209000000000000015500000000000000fb337c391c",
    x"030b0000000000000155fffffffffffff50003e5e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd8e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2eab1c",
    x"070a0000000000000155fffffffffffff8ef35ffa21c",
    x"08020000000000000155fffffffffffff6f669e7441c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7ac1c",
    x"0209000000000000015500000000000000fb337c331c",
    x"030b0000000000000155fffffffffffff50003e5ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd8b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ea51c",
    x"070a0000000000000155fffffffffffff8ef35ff9e1c",
    x"08020000000000000155fffffffffffff6f669e7421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7ad1c",
    x"0209000000000000015500000000000000fb337c2e1c",
    x"030b0000000000000155fffffffffffff50003e5eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43811c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e9f1c",
    x"070a0000000000000155fffffffffffff8ef35ff9b1c",
    x"08020000000000000155fffffffffffff6f669e73f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da0d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7af1c",
    x"0209000000000000015500000000000000fb337c281c",
    x"030b0000000000000155fffffffffffff50003e5ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f437d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e991c",
    x"070a0000000000000155fffffffffffff8ef35ff971c",
    x"08020000000000000155fffffffffffff6f669e73d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7b01c",
    x"0209000000000000015500000000000000fb337c231c",
    x"030b0000000000000155fffffffffffff50003e5ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e931c",
    x"070a0000000000000155fffffffffffff8ef35ff941c",
    x"08020000000000000155fffffffffffff6f669e73b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7b11c",
    x"0209000000000000015500000000000000fb337c1d1c",
    x"030b0000000000000155fffffffffffff50003e5ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e8d1c",
    x"070a0000000000000155fffffffffffff8ef35ff901c",
    x"08020000000000000155fffffffffffff6f669e7381c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266da011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7b21c",
    x"0209000000000000015500000000000000fb337c171c",
    x"030b0000000000000155fffffffffffff50003e5ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd7f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e861c",
    x"070a0000000000000155fffffffffffff8ef35ff8c1c",
    x"08020000000000000155fffffffffffff6f669e7361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d9fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7b31c",
    x"0209000000000000015500000000000000fb337c121c",
    x"030b0000000000000155fffffffffffff50003e5f01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd7d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f436e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e801c",
    x"070a0000000000000155fffffffffffff8ef35ff891c",
    x"08020000000000000155fffffffffffff6f669e7341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d9f81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe7b41c",
    x"0209000000000000025500000000000000fb337c0c1c",
    x"030b0000000000000255fffffffffffff50003e5f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dcd7b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f436b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2e7a1c",
    x"070a0000000000000255fffffffffffff8ef35ff851c",
    x"08020000000000000255fffffffffffff6f669e7311c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d9f41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7b51c",
    x"0209000000000000015500000000000000fb337c071c",
    x"030b0000000000000155fffffffffffff50003e5f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f43671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2e741c",
    x"070a0000000000000155fffffffffffff8ef35ff821c",
    x"08020000000000000155fffffffffffff6f669e72f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d9f01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7b61c",
    x"0209000000000000031f00000000000000fb337c011c",
    x"030b000000000000031ffffffffffffff50003e5f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcd761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f43631c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2e6e1c",
    x"070a000000000000031ffffffffffffff8ef35ff7e1c",
    x"0802000000000000031ffffffffffffff6f669e72c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d9ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7b71c",
    x"020900000000000000ae00000000000000fb337bfb1c",
    x"030b00000000000000aefffffffffffff50003e5f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcd731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f435f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2e681c",
    x"070a00000000000000aefffffffffffff8ef35ff7a1c",
    x"080200000000000000aefffffffffffff6f669e72a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d9e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7b81c",
    x"020900000000000001a400000000000000fb337bf61c",
    x"030b00000000000001a4fffffffffffff50003e5f51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcd711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f435c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2e621c",
    x"070a00000000000001a4fffffffffffff8ef35ff771c",
    x"080200000000000001a4fffffffffffff6f669e7281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d9e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe7ba1c",
    x"0209000000000000026600000000000000fb337bf01c",
    x"030b0000000000000266fffffffffffff50003e5f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dcd6f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f43581c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000266ffffffffffffff04cd2e5b1c",
    x"070a0000000000000266fffffffffffff8ef35ff731c",
    x"08020000000000000266fffffffffffff6f669e7251c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9df1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7bb1c",
    x"020900000000000002aa00000000000000fb337beb1c",
    x"030b00000000000002aafffffffffffff50003e5f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd6c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e551c",
    x"070a00000000000002aafffffffffffff8ef35ff701c",
    x"080200000000000002aafffffffffffff6f669e7231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9db1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7bc1c",
    x"020900000000000002aa00000000000000fb337be51c",
    x"030b00000000000002aafffffffffffff50003e5f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd6a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43511c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e4f1c",
    x"070a00000000000002aafffffffffffff8ef35ff6c1c",
    x"080200000000000002aafffffffffffff6f669e7201c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9d71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7bd1c",
    x"020900000000000002aa00000000000000fb337bdf1c",
    x"030b00000000000002aafffffffffffff50003e5f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f434d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e491c",
    x"070a00000000000002aafffffffffffff8ef35ff681c",
    x"080200000000000002aafffffffffffff6f669e71e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7be1c",
    x"020900000000000002aa00000000000000fb337bda1c",
    x"030b00000000000002aafffffffffffff50003e5fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e431c",
    x"070a00000000000002aafffffffffffff8ef35ff651c",
    x"080200000000000002aafffffffffffff6f669e71c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7bf1c",
    x"020900000000000002aa00000000000000fb337bd41c",
    x"030b00000000000002aafffffffffffff50003e5fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd631c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43461c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e3d1c",
    x"070a00000000000002aafffffffffffff8ef35ff611c",
    x"080200000000000002aafffffffffffff6f669e7191c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9ca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c01c",
    x"020900000000000002aa00000000000000fb337bcf1c",
    x"030b00000000000002aafffffffffffff50003e5fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e371c",
    x"070a00000000000002aafffffffffffff8ef35ff5e1c",
    x"080200000000000002aafffffffffffff6f669e7171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9c61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c11c",
    x"020900000000000002aa00000000000000fb337bc91c",
    x"030b00000000000002aafffffffffffff50003e5fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd5e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f433e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e301c",
    x"070a00000000000002aafffffffffffff8ef35ff5a1c",
    x"080200000000000002aafffffffffffff6f669e7151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9c21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c21c",
    x"020900000000000002aa00000000000000fb337bc31c",
    x"030b00000000000002aafffffffffffff50003e5fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd5b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f433a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e2a1c",
    x"070a00000000000002aafffffffffffff8ef35ff561c",
    x"080200000000000002aafffffffffffff6f669e7121c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c31c",
    x"020900000000000002aa00000000000000fb337bbe1c",
    x"030b00000000000002aafffffffffffff50003e5ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e241c",
    x"070a00000000000002aafffffffffffff8ef35ff531c",
    x"080200000000000002aafffffffffffff6f669e7101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c51c",
    x"020900000000000002aa00000000000000fb337bb81c",
    x"030b00000000000002aafffffffffffff50003e6001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43331c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e1e1c",
    x"070a00000000000002aafffffffffffff8ef35ff4f1c",
    x"080200000000000002aafffffffffffff6f669e70d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9b51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c61c",
    x"020900000000000002aa00000000000000fb337bb31c",
    x"030b00000000000002aafffffffffffff50003e6011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f432f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e181c",
    x"070a00000000000002aafffffffffffff8ef35ff4c1c",
    x"080200000000000002aafffffffffffff6f669e70b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9b11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c71c",
    x"020900000000000002aa00000000000000fb337bad1c",
    x"030b00000000000002aafffffffffffff50003e6021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f432c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e121c",
    x"070a00000000000002aafffffffffffff8ef35ff481c",
    x"080200000000000002aafffffffffffff6f669e7091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9ad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c81c",
    x"020900000000000002aa00000000000000fb337ba71c",
    x"030b00000000000002aafffffffffffff50003e6031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd4f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e0c1c",
    x"070a00000000000002aafffffffffffff8ef35ff441c",
    x"080200000000000002aafffffffffffff6f669e7061c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9a91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7c91c",
    x"020900000000000002aa00000000000000fb337ba21c",
    x"030b00000000000002aafffffffffffff50003e6041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd4d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2e051c",
    x"070a00000000000002aafffffffffffff8ef35ff411c",
    x"080200000000000002aafffffffffffff6f669e7041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7ca1c",
    x"020900000000000002aa00000000000000fb337b9c1c",
    x"030b00000000000002aafffffffffffff50003e6051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd4b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f43211c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2dff1c",
    x"070a00000000000002aafffffffffffff8ef35ff3d1c",
    x"080200000000000002aafffffffffffff6f669e7021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d9a01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7cb1c",
    x"020900000000000002aa00000000000000fb337b971c",
    x"030b00000000000002aafffffffffffff50003e6061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f431d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2df91c",
    x"070a00000000000002aafffffffffffff8ef35ff3a1c",
    x"080200000000000002aafffffffffffff6f669e6ff1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d99c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7cc1c",
    x"0209000000000000031f00000000000000fb337b911c",
    x"030b000000000000031ffffffffffffff50003e6071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcd461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f43191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2df31c",
    x"070a000000000000031ffffffffffffff8ef35ff361c",
    x"0802000000000000031ffffffffffffff6f669e6fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d9981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7cd1c",
    x"020900000000000000ae00000000000000fb337b8c1c",
    x"030b00000000000000aefffffffffffff50003e6081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcd431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f43161c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2ded1c",
    x"070a00000000000000aefffffffffffff8ef35ff321c",
    x"080200000000000000aefffffffffffff6f669e6fa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d9941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7ce1c",
    x"020900000000000001a400000000000000fb337b861c",
    x"030b00000000000001a4fffffffffffff50003e6091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcd411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f43121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2de71c",
    x"070a00000000000001a4fffffffffffff8ef35ff2f1c",
    x"080200000000000001a4fffffffffffff6f669e6f81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d9901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbe7d01c",
    x"020900000000000001aa00000000000000fb337b801c",
    x"030b00000000000001aafffffffffffff50003e60a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcd3f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f430e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd2de11c",
    x"070a00000000000001aafffffffffffff8ef35ff2b1c",
    x"080200000000000001aafffffffffffff6f669e6f61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d98b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe7d11c",
    x"0209000000000000029500000000000000fb337b7b1c",
    x"030b0000000000000295fffffffffffff50003e60b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcd3c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f430a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2dda1c",
    x"070a0000000000000295fffffffffffff8ef35ff281c",
    x"08020000000000000295fffffffffffff6f669e6f31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266d9871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe7d21c",
    x"0209000000000000015a00000000000000fb337b751c",
    x"030b000000000000015afffffffffffff50003e60c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dcd3a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f43071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd2dd41c",
    x"070a000000000000015afffffffffffff8ef35ff241c",
    x"0802000000000000015afffffffffffff6f669e6f11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d9831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe7d31c",
    x"0209000000000000025500000000000000fb337b701c",
    x"030b0000000000000255fffffffffffff50003e60d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dcd371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f43031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2dce1c",
    x"070a0000000000000255fffffffffffff8ef35ff201c",
    x"08020000000000000255fffffffffffff6f669e6ee1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d97f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe7d41c",
    x"0209000000000000015600000000000000fb337b6a1c",
    x"030b00000000000002aafffffffffffff50003e60e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcd351c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f42ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd2dc81c",
    x"070a00000000000002aafffffffffffff8ef35ff1d1c",
    x"08020000000000000156fffffffffffff6f669e6ec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d97b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7d51c",
    x"0209000000000000016500000000000000fb337b641c",
    x"030b000000000000019afffffffffffff50003e60f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcd331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a90000000000000b072f42fc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd2dc21c",
    x"070a00000000000001aafffffffffffff8ef35ff191c",
    x"08020000000000000156fffffffffffff6f669e6ea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d9771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe7d61c",
    x"020900000000000002a500000000000000fb337b5f1c",
    x"030b000000000000019afffffffffffff50003e6101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcd301c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd2dbc1c",
    x"070a0000000000000165fffffffffffff8ef35ff161c",
    x"08020000000000000265fffffffffffff6f669e6e71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d9721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe7d71c",
    x"0209000000000000026600000000000000fb337b591c",
    x"030b0000000000000299fffffffffffff50003e6111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dcd2e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f42f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2db61c",
    x"070a0000000000000256fffffffffffff8ef35ff121c",
    x"08020000000000000195fffffffffffff6f669e6e51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266d96e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe7d81c",
    x"0209000000000000029900000000000000fb337b541c",
    x"030b0000000000000259fffffffffffff50003e6121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcd2b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f42f11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd2daf1c",
    x"070a0000000000000266fffffffffffff8ef35ff0e1c",
    x"080200000000000001a5fffffffffffff6f669e6e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266d96a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7d91c",
    x"020900000000000002aa00000000000000fb337b4e1c",
    x"030b00000000000002a5fffffffffffff50003e6131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dcd291c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f42ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd2da91c",
    x"070a0000000000000295fffffffffffff8ef35ff0b1c",
    x"080200000000000001a5fffffffffffff6f669e6e01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266d9661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe7db1c",
    x"020900000000000002a500000000000000fb337b481c",
    x"030b000000000000016afffffffffffff50003e6141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f42e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd2da31c",
    x"070a0000000000000255fffffffffffff8ef35ff071c",
    x"08020000000000000169fffffffffffff6f669e6de1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266d9621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe7dc1c",
    x"0209000000000000025600000000000000fb337b431c",
    x"030b0000000000000166fffffffffffff50003e6151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcd241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f42e61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2d9d1c",
    x"070a000000000000029afffffffffffff8ef35ff041c",
    x"08020000000000000295fffffffffffff6f669e6db1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000269ffffffffffffff0266d95d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbe7dd1c",
    x"0209000000000000015500000000000000fb337b3d1c",
    x"030b0000000000000296fffffffffffff50003e6161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dcd221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f42e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd2d971c",
    x"070a0000000000000156fffffffffffff8ef35ff001c",
    x"08020000000000000266fffffffffffff6f669e6d91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d9591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe7de1c",
    x"0209000000000000016500000000000000fb337b381c",
    x"030b0000000000000265fffffffffffff50003e6171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dcd1f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f42de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000265ffffffffffffff04cd2d911c",
    x"070a0000000000000295fffffffffffff8ef35fefc1c",
    x"0802000000000000029afffffffffffff6f669e6d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d9551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a90000000000000b0bfbe7df1c",
    x"0209000000000000015900000000000000fb337b321c",
    x"030b00000000000002a5fffffffffffff50003e6181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dcd1d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f42da1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd2d8b1c",
    x"070a00000000000001a5fffffffffffff8ef35fef91c",
    x"080200000000000001a5fffffffffffff6f669e6d41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d9511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbe7e01c",
    x"0209000000000000016500000000000000fb337b2c1c",
    x"030b00000000000001aafffffffffffff50003e6191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd1b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f42d71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2d841c",
    x"070a0000000000000296fffffffffffff8ef35fef51c",
    x"08020000000000000266fffffffffffff6f669e6d21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266d94d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7e11c",
    x"0209000000000000015a00000000000000fb337b271c",
    x"030b00000000000002a5fffffffffffff50003e61a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dcd181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f42d31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2d7e1c",
    x"070a00000000000002a5fffffffffffff8ef35fef21c",
    x"08020000000000000169fffffffffffff6f669e6cf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d9481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7e21c",
    x"0209000000000000031f00000000000000fb337b211c",
    x"030b000000000000031ffffffffffffff50003e61b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcd161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f42cf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2d781c",
    x"070a000000000000031ffffffffffffff8ef35feee1c",
    x"0802000000000000031ffffffffffffff6f669e6cd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d9441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7e31c",
    x"020900000000000000ae00000000000000fb337b1c1c",
    x"030b00000000000000aefffffffffffff50003e61c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcd131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f42cc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2d721c",
    x"070a00000000000000aefffffffffffff8ef35feea1c",
    x"080200000000000000aefffffffffffff6f669e6cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d9401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7e51c",
    x"020900000000000001a400000000000000fb337b161c",
    x"030b00000000000001a4fffffffffffff50003e61d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcd111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f42c81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2d6c1c",
    x"070a00000000000001a4fffffffffffff8ef35fee71c",
    x"080200000000000001a4fffffffffffff6f669e6c81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d93c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe7e61c",
    x"0209000000000000016a00000000000000fb337b101c",
    x"030b000000000000016afffffffffffff50003e61e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcd0f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f42c41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd2d661c",
    x"070a000000000000016afffffffffffff8ef35fee31c",
    x"0802000000000000016afffffffffffff6f669e6c61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d9381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7e71c",
    x"0209000000000000015500000000000000fb337b0b1c",
    x"030b0000000000000155fffffffffffff50003e61f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcd0c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42c11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2d5f1c",
    x"070a0000000000000155fffffffffffff8ef35fee01c",
    x"08020000000000000155fffffffffffff6f669e6c31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266d9331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe7e81c",
    x"0209000000000000019500000000000000fb337b051c",
    x"030b0000000000000195fffffffffffff50003e6201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dcd0a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f42bd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2d591c",
    x"070a0000000000000195fffffffffffff8ef35fedc1c",
    x"080200000000000002a5fffffffffffff6f669e6c11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d92f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7e91c",
    x"020900000000000002aa00000000000000fb337b001c",
    x"030b00000000000002aafffffffffffff50003e6211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcd071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f42b91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2d531c",
    x"070a00000000000002aafffffffffffff8ef35fed81c",
    x"08020000000000000155fffffffffffff6f669e6bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d92b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe7ea1c",
    x"0209000000000000029600000000000000fb337afa1c",
    x"030b00000000000001aafffffffffffff50003e6221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dcd051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f42b61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2d4d1c",
    x"070a0000000000000256fffffffffffff8ef35fed51c",
    x"08020000000000000155fffffffffffff6f669e6bc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266d9271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe7eb1c",
    x"0209000000000000026500000000000000fb337af41c",
    x"030b00000000000002a9fffffffffffff50003e6231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dcd031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f42b21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd2d471c",
    x"070a000000000000029afffffffffffff8ef35fed11c",
    x"08020000000000000159fffffffffffff6f669e6ba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266d9231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe7ec1c",
    x"0209000000000000029600000000000000fb337aef1c",
    x"030b000000000000016afffffffffffff50003e6241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dcd001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f42ae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd2d411c",
    x"070a0000000000000159fffffffffffff8ef35fecd1c",
    x"0802000000000000015afffffffffffff6f669e6b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d91e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe7ed1c",
    x"0209000000000000016900000000000000fb337ae91c",
    x"030b0000000000000295fffffffffffff50003e6251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dccfe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f42aa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd2d3b1c",
    x"070a0000000000000196fffffffffffff8ef35feca1c",
    x"08020000000000000299fffffffffffff6f669e6b51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d91a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe7ee1c",
    x"020900000000000002a500000000000000fb337ae41c",
    x"030b0000000000000156fffffffffffff50003e6261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dccfb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f42a71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd2d341c",
    x"070a00000000000002a6fffffffffffff8ef35fec61c",
    x"080200000000000001a5fffffffffffff6f669e6b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266d9161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe7f01c",
    x"0209000000000000025500000000000000fb337ade1c",
    x"030b000000000000016afffffffffffff50003e6271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dccf91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f42a31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2d2e1c",
    x"070a0000000000000295fffffffffffff8ef35fec31c",
    x"0802000000000000026afffffffffffff6f669e6b01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d9121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe7f11c",
    x"0209000000000000029a00000000000000fb337ad81c",
    x"030b0000000000000269fffffffffffff50003e6281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dccf71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f429f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2d281c",
    x"070a0000000000000196fffffffffffff8ef35febf1c",
    x"08020000000000000165fffffffffffff6f669e6ae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d90e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe7f21c",
    x"020900000000000001a600000000000000fb337ad31c",
    x"030b000000000000019afffffffffffff50003e6291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dccf41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f429c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd2d221c",
    x"070a000000000000026afffffffffffff8ef35febb1c",
    x"0802000000000000019afffffffffffff6f669e6ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266d90a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbe7f31c",
    x"0209000000000000025a00000000000000fb337acd1c",
    x"030b00000000000002a9fffffffffffff50003e62a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dccf21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f42981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd2d1c1c",
    x"070a00000000000002a6fffffffffffff8ef35feb81c",
    x"08020000000000000295fffffffffffff6f669e6a91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d9051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe7f41c",
    x"0209000000000000029600000000000000fb337ac81c",
    x"030b000000000000025afffffffffffff50003e62b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dccef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f42941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd2d161c",
    x"070a000000000000019afffffffffffff8ef35feb41c",
    x"0802000000000000029afffffffffffff6f669e6a71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266d9011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe7f51c",
    x"0209000000000000019900000000000000fb337ac21c",
    x"030b0000000000000156fffffffffffff50003e62c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcced1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f42911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd2d101c",
    x"070a0000000000000166fffffffffffff8ef35feb11c",
    x"080200000000000001a9fffffffffffff6f669e6a41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d8fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe7f61c",
    x"0209000000000000015600000000000000fb337abc1c",
    x"030b0000000000000169fffffffffffff50003e62d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dcceb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f428d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd2d091c",
    x"070a0000000000000159fffffffffffff8ef35fead1c",
    x"08020000000000000255fffffffffffff6f669e6a21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266d8f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7f71c",
    x"0209000000000000029a00000000000000fb337ab71c",
    x"030b00000000000002a9fffffffffffff50003e62e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcce81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd2d031c",
    x"070a0000000000000159fffffffffffff8ef35fea91c",
    x"08020000000000000299fffffffffffff6f669e6a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d8f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe7f81c",
    x"0209000000000000031f00000000000000fb337ab11c",
    x"030b000000000000031ffffffffffffff50003e62f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcce61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f42861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2cfd1c",
    x"070a000000000000031ffffffffffffff8ef35fea61c",
    x"0802000000000000031ffffffffffffff6f669e69d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d8f01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe7f91c",
    x"020900000000000000ae00000000000000fb337aac1c",
    x"030b00000000000000aefffffffffffff50003e6301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcce31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f42821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2cf71c",
    x"070a00000000000000aefffffffffffff8ef35fea21c",
    x"080200000000000000aefffffffffffff6f669e69b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d8ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe7fb1c",
    x"020900000000000001a400000000000000fb337aa61c",
    x"030b00000000000001a4fffffffffffff50003e6311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcce11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f427e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2cf11c",
    x"070a00000000000001a4fffffffffffff8ef35fe9f1c",
    x"080200000000000001a4fffffffffffff6f669e6991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266d8e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe7fc1c",
    x"0209000000000000026a00000000000000fb337aa01c",
    x"030b000000000000026afffffffffffff50003e6321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dccdf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f427a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026affffffffffffff04cd2ceb1c",
    x"070a000000000000026afffffffffffff8ef35fe9b1c",
    x"0802000000000000026afffffffffffff6f669e6961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7fd1c",
    x"0209000000000000015500000000000000fb337a9b1c",
    x"030b0000000000000155fffffffffffff50003e6331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dccdc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f42771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd2ce51c",
    x"070a00000000000002a9fffffffffffff8ef35fe971c",
    x"08020000000000000155fffffffffffff6f669e6941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe7fe1c",
    x"0209000000000000015500000000000000fb337a951c",
    x"030b0000000000000155fffffffffffff50003e6341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dccda1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f42731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2cde1c",
    x"070a00000000000001aafffffffffffff8ef35fe941c",
    x"08020000000000000155fffffffffffff6f669e6911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266d8db1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe7ff1c",
    x"0209000000000000015600000000000000fb337a901c",
    x"030b0000000000000155fffffffffffff50003e6351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dccd71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f426f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd2cd81c",
    x"070a00000000000002aafffffffffffff8ef35fe901c",
    x"08020000000000000155fffffffffffff6f669e68f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d8d71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe8001c",
    x"0209000000000000025500000000000000fb337a8a1c",
    x"030b0000000000000195fffffffffffff50003e6361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dccd51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f426c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd2cd21c",
    x"070a000000000000026afffffffffffff8ef35fe8d1c",
    x"08020000000000000195fffffffffffff6f669e68d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d8d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe8011c",
    x"0209000000000000016500000000000000fb337a841c",
    x"030b00000000000002a9fffffffffffff50003e6371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dccd21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000259ffffffffffffff04cd2ccc1c",
    x"070a0000000000000256fffffffffffff8ef35fe891c",
    x"08020000000000000299fffffffffffff6f669e68a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d8cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe8021c",
    x"0209000000000000019900000000000000fb337a7f1c",
    x"030b0000000000000195fffffffffffff50003e6381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dccd01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f42641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd2cc61c",
    x"070a0000000000000266fffffffffffff8ef35fe851c",
    x"080200000000000002a6fffffffffffff6f669e6881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d8cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe8031c",
    x"0209000000000000016500000000000000fb337a791c",
    x"030b0000000000000166fffffffffffff50003e6391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dccce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f42611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd2cc01c",
    x"070a0000000000000156fffffffffffff8ef35fe821c",
    x"0802000000000000025afffffffffffff6f669e6851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d8c61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe8041c",
    x"0209000000000000019500000000000000fb337a741c",
    x"030b0000000000000265fffffffffffff50003e63a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dcccb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f425d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd2cba1c",
    x"070a000000000000025afffffffffffff8ef35fe7e1c",
    x"0802000000000000016afffffffffffff6f669e6831c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d8c21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe8061c",
    x"0209000000000000026a00000000000000fb337a6e1c",
    x"030b00000000000002aafffffffffffff50003e63b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dccc91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f42591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd2cb31c",
    x"070a0000000000000195fffffffffffff8ef35fe7b1c",
    x"08020000000000000195fffffffffffff6f669e6811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266d8be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe8071c",
    x"0209000000000000025600000000000000fb337a681c",
    x"030b00000000000002a5fffffffffffff50003e63c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dccc61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f42561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd2cad1c",
    x"070a00000000000002a5fffffffffffff8ef35fe771c",
    x"08020000000000000295fffffffffffff6f669e67e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d8ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe8081c",
    x"020900000000000001a900000000000000fb337a631c",
    x"030b0000000000000155fffffffffffff50003e63d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dccc41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f42521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd2ca71c",
    x"070a0000000000000256fffffffffffff8ef35fe731c",
    x"08020000000000000199fffffffffffff6f669e67c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d8b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe8091c",
    x"0209000000000000029500000000000000fb337a5d1c",
    x"030b0000000000000299fffffffffffff50003e63e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dccc21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f424e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd2ca11c",
    x"070a0000000000000266fffffffffffff8ef35fe701c",
    x"08020000000000000166fffffffffffff6f669e67a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d8b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe80a1c",
    x"0209000000000000016900000000000000fb337a581c",
    x"030b000000000000016afffffffffffff50003e63f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dccbf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f424a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd2c9b1c",
    x"070a0000000000000256fffffffffffff8ef35fe6c1c",
    x"08020000000000000199fffffffffffff6f669e6771c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266d8ad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe80b1c",
    x"0209000000000000026a00000000000000fb337a521c",
    x"030b000000000000016afffffffffffff50003e6401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dccbd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f42471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd2c951c",
    x"070a00000000000001a5fffffffffffff8ef35fe681c",
    x"08020000000000000266fffffffffffff6f669e6751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d8a91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe80c1c",
    x"020900000000000001a900000000000000fb337a4c1c",
    x"030b000000000000026afffffffffffff50003e6411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dccba1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f42431c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd2c8e1c",
    x"070a0000000000000166fffffffffffff8ef35fe651c",
    x"08020000000000000296fffffffffffff6f669e6721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266d8a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe80d1c",
    x"020900000000000002a600000000000000fb337a471c",
    x"030b000000000000015afffffffffffff50003e6421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dccb81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f423f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd2c881c",
    x"070a0000000000000295fffffffffffff8ef35fe611c",
    x"080200000000000002a5fffffffffffff6f669e6701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d8a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe80e1c",
    x"0209000000000000031f00000000000000fb337a411c",
    x"030b000000000000031ffffffffffffff50003e6431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dccb61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f423c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2c821c",
    x"070a000000000000031ffffffffffffff8ef35fe5e1c",
    x"0802000000000000031ffffffffffffff6f669e66e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d89d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8101c",
    x"020900000000000000ae00000000000000fb337a3c1c",
    x"030b00000000000000aefffffffffffff50003e6441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dccb31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f42381c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2c7c1c",
    x"070a00000000000000aefffffffffffff8ef35fe5a1c",
    x"080200000000000000aefffffffffffff6f669e66b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d8981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8111c",
    x"020900000000000001a400000000000000fb337a361c",
    x"030b00000000000001a4fffffffffffff50003e6451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dccb11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f42341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2c761c",
    x"070a00000000000001a4fffffffffffff8ef35fe561c",
    x"080200000000000001a4fffffffffffff6f669e6691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266d8941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe8121c",
    x"0209000000000000015a00000000000000fb337a301c",
    x"030b000000000000015afffffffffffff50003e6461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dccae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f42311c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd2c701c",
    x"070a000000000000015afffffffffffff8ef35fe531c",
    x"0802000000000000015afffffffffffff6f669e6661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d8901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8131c",
    x"020900000000000001aa00000000000000fb337a2b1c",
    x"030b0000000000000255fffffffffffff50003e6471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dccac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f422d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2c6a1c",
    x"070a0000000000000155fffffffffffff8ef35fe4f1c",
    x"08020000000000000155fffffffffffff6f669e6641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266d88c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe8141c",
    x"0209000000000000016900000000000000fb337a251c",
    x"030b0000000000000269fffffffffffff50003e6481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dccaa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f42291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd2c631c",
    x"070a00000000000002a6fffffffffffff8ef35fe4c1c",
    x"080200000000000001a5fffffffffffff6f669e6621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266d8881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe8151c",
    x"020900000000000001a600000000000000fb337a201c",
    x"030b0000000000000296fffffffffffff50003e6491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dcca71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f42261c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd2c5d1c",
    x"070a000000000000029afffffffffffff8ef35fe481c",
    x"08020000000000000196fffffffffffff6f669e65f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d8831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe8161c",
    x"0209000000000000026900000000000000fb337a1a1c",
    x"030b0000000000000255fffffffffffff50003e64a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dcca51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f42221c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000199ffffffffffffff04cd2c571c",
    x"070a0000000000000265fffffffffffff8ef35fe441c",
    x"08020000000000000256fffffffffffff6f669e65d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d87f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe8171c",
    x"0209000000000000015600000000000000fb337a141c",
    x"030b0000000000000155fffffffffffff50003e64b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcca21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f421e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd2c511c",
    x"070a00000000000002aafffffffffffff8ef35fe411c",
    x"08020000000000000155fffffffffffff6f669e65b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d87b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8181c",
    x"0209000000000000015500000000000000fb337a0f1c",
    x"030b0000000000000155fffffffffffff50003e64c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcca01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f421a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2c4b1c",
    x"070a00000000000002aafffffffffffff8ef35fe3d1c",
    x"08020000000000000155fffffffffffff6f669e6581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8191c",
    x"020900000000000002aa00000000000000fb337a091c",
    x"030b00000000000002aafffffffffffff50003e64d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc9e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2c451c",
    x"070a0000000000000155fffffffffffff8ef35fe3a1c",
    x"080200000000000002aafffffffffffff6f669e6561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe81b1c",
    x"020900000000000002aa00000000000000fb337a041c",
    x"030b00000000000002aafffffffffffff50003e64e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc9b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42131c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2c3f1c",
    x"070a0000000000000155fffffffffffff8ef35fe361c",
    x"080200000000000002aafffffffffffff6f669e6531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d86e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe81c1c",
    x"020900000000000002aa00000000000000fb3379fe1c",
    x"030b00000000000002aafffffffffffff50003e64f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc991c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f420f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2c381c",
    x"070a0000000000000155fffffffffffff8ef35fe321c",
    x"080200000000000002aafffffffffffff6f669e6511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266d86a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbe81d1c",
    x"020900000000000001a600000000000000fb3379f81c",
    x"030b00000000000001a6fffffffffffff50003e6501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000259fffffffffffff4099dcc961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f420c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd2c321c",
    x"070a0000000000000259fffffffffffff8ef35fe2f1c",
    x"080200000000000001a6fffffffffffff6f669e64f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe81e1c",
    x"020900000000000002aa00000000000000fb3379f31c",
    x"030b00000000000002aafffffffffffff50003e6511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc941c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42081c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2c2c1c",
    x"070a0000000000000155fffffffffffff8ef35fe2b1c",
    x"080200000000000002aafffffffffffff6f669e64c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe81f1c",
    x"020900000000000002aa00000000000000fb3379ed1c",
    x"030b00000000000002aafffffffffffff50003e6521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc921c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f42041c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2c261c",
    x"070a0000000000000155fffffffffffff8ef35fe271c",
    x"080200000000000002aafffffffffffff6f669e64a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d85e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe8201c",
    x"020900000000000002a600000000000000fb3379e81c",
    x"030b00000000000002a6fffffffffffff50003e6531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcc8f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f42011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd2c201c",
    x"070a0000000000000159fffffffffffff8ef35fe241c",
    x"080200000000000002a6fffffffffffff6f669e6471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d85a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a50000000000000b0bfbe8211c",
    x"0209000000000000029500000000000000fb3379e21c",
    x"030b00000000000002aafffffffffffff50003e6541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dcc8d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f41fd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd2c1a1c",
    x"070a000000000000019afffffffffffff8ef35fe201c",
    x"080200000000000002a5fffffffffffff6f669e6451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d8551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe8221c",
    x"0209000000000000016a00000000000000fb3379dd1c",
    x"030b000000000000016afffffffffffff50003e6551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcc8a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002650000000000000b072f41f91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd2c141c",
    x"070a0000000000000265fffffffffffff8ef35fe1d1c",
    x"080200000000000001aafffffffffffff6f669e6431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d8511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe8231c",
    x"0209000000000000015a00000000000000fb3379d71c",
    x"030b000000000000015afffffffffffff50003e6561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dcc881c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f41f61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd2c0d1c",
    x"070a00000000000002a5fffffffffffff8ef35fe191c",
    x"0802000000000000015afffffffffffff6f669e6401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d84d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8251c",
    x"0209000000000000031f00000000000000fb3379d11c",
    x"030b000000000000031ffffffffffffff50003e6571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcc851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f41f21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2c071c",
    x"070a000000000000031ffffffffffffff8ef35fe151c",
    x"0802000000000000031ffffffffffffff6f669e63e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d8491c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8261c",
    x"020900000000000000ae00000000000000fb3379cc1c",
    x"030b00000000000000aefffffffffffff50003e6581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcc831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f41ee1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2c011c",
    x"070a00000000000000aefffffffffffff8ef35fe121c",
    x"080200000000000000aefffffffffffff6f669e63b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d8451c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8271c",
    x"020900000000000001a400000000000000fb3379c61c",
    x"030b00000000000001a4fffffffffffff50003e6591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcc811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f41eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2bfb1c",
    x"070a00000000000001a4fffffffffffff8ef35fe0e1c",
    x"080200000000000001a4fffffffffffff6f669e6391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266d8401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe8281c",
    x"0209000000000000025a00000000000000fb3379c11c",
    x"030b000000000000025afffffffffffff50003e65a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dcc7e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f41e71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd2bf51c",
    x"070a000000000000025afffffffffffff8ef35fe0b1c",
    x"0802000000000000025afffffffffffff6f669e6371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d83c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8291c",
    x"020900000000000002aa00000000000000fb3379bb1c",
    x"030b00000000000002aafffffffffffff50003e65b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc7c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41e31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bef1c",
    x"070a00000000000002aafffffffffffff8ef35fe071c",
    x"080200000000000002aafffffffffffff6f669e6341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d8381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe82a1c",
    x"0209000000000000029a00000000000000fb3379b51c",
    x"030b000000000000029afffffffffffff50003e65c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcc791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f41df1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd2be81c",
    x"070a000000000000029afffffffffffff8ef35fe031c",
    x"0802000000000000029afffffffffffff6f669e6321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d8341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe82b1c",
    x"020900000000000002aa00000000000000fb3379b01c",
    x"030b00000000000002aafffffffffffff50003e65d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41dc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2be21c",
    x"070a00000000000002aafffffffffffff8ef35fe001c",
    x"080200000000000002aafffffffffffff6f669e6301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d8301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe82c1c",
    x"020900000000000002aa00000000000000fb3379aa1c",
    x"030b00000000000002aafffffffffffff50003e65e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41d81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bdc1c",
    x"070a00000000000002aafffffffffffff8ef35fdfc1c",
    x"080200000000000002aafffffffffffff6f669e62d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d82b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe82d1c",
    x"020900000000000002aa00000000000000fb3379a51c",
    x"030b00000000000002aafffffffffffff50003e65f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc721c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41d41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bd61c",
    x"070a00000000000002aafffffffffffff8ef35fdf91c",
    x"080200000000000002aafffffffffffff6f669e62b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d8271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe82e1c",
    x"020900000000000002aa00000000000000fb33799f1c",
    x"030b00000000000002aafffffffffffff50003e6601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bd01c",
    x"070a00000000000002aafffffffffffff8ef35fdf51c",
    x"080200000000000002aafffffffffffff6f669e6281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d8231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8301c",
    x"020900000000000002aa00000000000000fb3379991c",
    x"030b00000000000002aafffffffffffff50003e6611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc6d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41cd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bca1c",
    x"070a00000000000002aafffffffffffff8ef35fdf11c",
    x"080200000000000002aafffffffffffff6f669e6261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d81f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8311c",
    x"020900000000000002aa00000000000000fb3379941c",
    x"030b00000000000002aafffffffffffff50003e6621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc6b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bc41c",
    x"070a00000000000002aafffffffffffff8ef35fdee1c",
    x"080200000000000002aafffffffffffff6f669e6241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d81b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8321c",
    x"020900000000000002aa00000000000000fb33798e1c",
    x"030b00000000000002aafffffffffffff50003e6631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41c61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2bbd1c",
    x"070a00000000000002aafffffffffffff8ef35fdea1c",
    x"080200000000000002aafffffffffffff6f669e6211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d8161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe8331c",
    x"0209000000000000016600000000000000fb3379891c",
    x"030b0000000000000166fffffffffffff50003e6641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dcc661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f41c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd2bb71c",
    x"070a0000000000000166fffffffffffff8ef35fde61c",
    x"08020000000000000166fffffffffffff6f669e61f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8341c",
    x"0209000000000000015500000000000000fb3379831c",
    x"030b0000000000000155fffffffffffff50003e6651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2bb11c",
    x"070a0000000000000155fffffffffffff8ef35fde31c",
    x"08020000000000000155fffffffffffff6f669e61c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d80e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8351c",
    x"0209000000000000015500000000000000fb33797d1c",
    x"030b0000000000000155fffffffffffff50003e6661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41bb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2bab1c",
    x"070a0000000000000155fffffffffffff8ef35fddf1c",
    x"08020000000000000155fffffffffffff6f669e61a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d80a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8361c",
    x"0209000000000000015500000000000000fb3379781c",
    x"030b0000000000000155fffffffffffff50003e6671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc5f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ba51c",
    x"070a0000000000000155fffffffffffff8ef35fddc1c",
    x"08020000000000000155fffffffffffff6f669e6181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8371c",
    x"0209000000000000015500000000000000fb3379721c",
    x"030b0000000000000155fffffffffffff50003e6681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc5d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2b9f1c",
    x"070a0000000000000155fffffffffffff8ef35fdd81c",
    x"08020000000000000155fffffffffffff6f669e6151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d8021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8381c",
    x"0209000000000000015500000000000000fb33796d1c",
    x"030b0000000000000155fffffffffffff50003e6681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc5a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2b991c",
    x"070a0000000000000155fffffffffffff8ef35fdd41c",
    x"08020000000000000155fffffffffffff6f669e6131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d7fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe83a1c",
    x"0209000000000000015900000000000000fb3379671c",
    x"030b0000000000000159fffffffffffff50003e6691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dcc581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f41ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd2b921c",
    x"070a0000000000000159fffffffffffff8ef35fdd11c",
    x"08020000000000000159fffffffffffff6f669e6111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d7f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe83b1c",
    x"0209000000000000031f00000000000000fb3379611c",
    x"030b000000000000031ffffffffffffff50003e66a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcc551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f41a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2b8c1c",
    x"070a000000000000031ffffffffffffff8ef35fdcd1c",
    x"0802000000000000031ffffffffffffff6f669e60e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d7f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe83c1c",
    x"020900000000000000ae00000000000000fb33795c1c",
    x"030b00000000000000aefffffffffffff50003e66b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcc531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f41a41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2b861c",
    x"070a00000000000000aefffffffffffff8ef35fdca1c",
    x"080200000000000000aefffffffffffff6f669e60c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d7f11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe83d1c",
    x"020900000000000001a400000000000000fb3379561c",
    x"030b00000000000001a4fffffffffffff50003e66c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcc501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f41a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2b801c",
    x"070a00000000000001a4fffffffffffff8ef35fdc61c",
    x"080200000000000001a4fffffffffffff6f669e6091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d7ed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe83e1c",
    x"0209000000000000029a00000000000000fb3379511c",
    x"030b000000000000029afffffffffffff50003e66d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcc4e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f419d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd2b7a1c",
    x"070a000000000000029afffffffffffff8ef35fdc21c",
    x"0802000000000000029afffffffffffff6f669e6071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe83f1c",
    x"020900000000000002aa00000000000000fb33794b1c",
    x"030b00000000000002aafffffffffffff50003e66e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc4c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41991c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b741c",
    x"070a00000000000002aafffffffffffff8ef35fdbf1c",
    x"080200000000000002aafffffffffffff6f669e6051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8401c",
    x"020900000000000002aa00000000000000fb3379451c",
    x"030b00000000000002aafffffffffffff50003e66f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b6e1c",
    x"070a00000000000002aafffffffffffff8ef35fdbb1c",
    x"080200000000000002aafffffffffffff6f669e6021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8411c",
    x"020900000000000002aa00000000000000fb3379401c",
    x"030b00000000000002aafffffffffffff50003e6701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b671c",
    x"070a00000000000002aafffffffffffff8ef35fdb71c",
    x"080200000000000002aafffffffffffff6f669e6001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7dc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8421c",
    x"020900000000000002aa00000000000000fb33793a1c",
    x"030b00000000000002aafffffffffffff50003e6711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f418e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b611c",
    x"070a00000000000002aafffffffffffff8ef35fdb41c",
    x"080200000000000002aafffffffffffff6f669e5fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8431c",
    x"020900000000000002aa00000000000000fb3379351c",
    x"030b00000000000002aafffffffffffff50003e6721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f418b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b5b1c",
    x"070a00000000000002aafffffffffffff8ef35fdb01c",
    x"080200000000000002aafffffffffffff6f669e5fb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8451c",
    x"020900000000000002aa00000000000000fb33792f1c",
    x"030b00000000000002aafffffffffffff50003e6731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc401c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b551c",
    x"070a00000000000002aafffffffffffff8ef35fdad1c",
    x"080200000000000002aafffffffffffff6f669e5f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8461c",
    x"020900000000000002aa00000000000000fb3379291c",
    x"030b00000000000002aafffffffffffff50003e6741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc3d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41831c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b4f1c",
    x"070a00000000000002aafffffffffffff8ef35fda91c",
    x"080200000000000002aafffffffffffff6f669e5f61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8471c",
    x"020900000000000002aa00000000000000fb3379241c",
    x"030b00000000000002aafffffffffffff50003e6751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc3b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b491c",
    x"070a00000000000002aafffffffffffff8ef35fda51c",
    x"080200000000000002aafffffffffffff6f669e5f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8481c",
    x"020900000000000002aa00000000000000fb33791e1c",
    x"030b00000000000002aafffffffffffff50003e6761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f417c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b421c",
    x"070a00000000000002aafffffffffffff8ef35fda21c",
    x"080200000000000002aafffffffffffff6f669e5f11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8491c",
    x"020900000000000002aa00000000000000fb3379191c",
    x"030b00000000000002aafffffffffffff50003e6771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b3c1c",
    x"070a00000000000002aafffffffffffff8ef35fd9e1c",
    x"080200000000000002aafffffffffffff6f669e5ef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe84a1c",
    x"020900000000000002aa00000000000000fb3379131c",
    x"030b00000000000002aafffffffffffff50003e6781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b361c",
    x"070a00000000000002aafffffffffffff8ef35fd9b1c",
    x"080200000000000002aafffffffffffff6f669e5ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe84b1c",
    x"020900000000000002aa00000000000000fb33790d1c",
    x"030b00000000000002aafffffffffffff50003e6791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b301c",
    x"070a00000000000002aafffffffffffff8ef35fd971c",
    x"080200000000000002aafffffffffffff6f669e5ea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe84c1c",
    x"020900000000000002aa00000000000000fb3379081c",
    x"030b00000000000002aafffffffffffff50003e67a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc2f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f416d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b2a1c",
    x"070a00000000000002aafffffffffffff8ef35fd931c",
    x"080200000000000002aafffffffffffff6f669e5e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe84d1c",
    x"020900000000000002aa00000000000000fb3379021c",
    x"030b00000000000002aafffffffffffff50003e67b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc2c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f416a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b241c",
    x"070a00000000000002aafffffffffffff8ef35fd901c",
    x"080200000000000002aafffffffffffff6f669e5e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d7ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe84f1c",
    x"0209000000000000029a00000000000000fb3378fd1c",
    x"030b000000000000029afffffffffffff50003e67c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcc2a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f41661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd2b1e1c",
    x"070a000000000000029afffffffffffff8ef35fd8c1c",
    x"0802000000000000029afffffffffffff6f669e5e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8501c",
    x"020900000000000002aa00000000000000fb3378f71c",
    x"030b00000000000002aafffffffffffff50003e67d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcc281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f41621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2b171c",
    x"070a00000000000002aafffffffffffff8ef35fd881c",
    x"080200000000000002aafffffffffffff6f669e5e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d7a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8511c",
    x"0209000000000000031f00000000000000fb3378f11c",
    x"030b000000000000031ffffffffffffff50003e67e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcc251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f415e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2b111c",
    x"070a000000000000031ffffffffffffff8ef35fd851c",
    x"0802000000000000031ffffffffffffff6f669e5de1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d7a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8521c",
    x"020900000000000000ae00000000000000fb3378ec1c",
    x"030b00000000000000aefffffffffffff50003e67f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcc231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f415b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2b0b1c",
    x"070a00000000000000aefffffffffffff8ef35fd811c",
    x"080200000000000000aefffffffffffff6f669e5dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d79d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8531c",
    x"020900000000000001a400000000000000fb3378e61c",
    x"030b00000000000001a4fffffffffffff50003e6801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcc201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f41571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2b051c",
    x"070a00000000000001a4fffffffffffff8ef35fd7e1c",
    x"080200000000000001a4fffffffffffff6f669e5da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266d7991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe8541c",
    x"0209000000000000019a00000000000000fb3378e11c",
    x"030b000000000000019afffffffffffff50003e6811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dcc1e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f41531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd2aff1c",
    x"070a000000000000019afffffffffffff8ef35fd7a1c",
    x"0802000000000000019afffffffffffff6f669e5d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8551c",
    x"0209000000000000015500000000000000fb3378db1c",
    x"030b0000000000000155fffffffffffff50003e6821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc1b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2af91c",
    x"070a0000000000000155fffffffffffff8ef35fd761c",
    x"08020000000000000155fffffffffffff6f669e5d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8561c",
    x"0209000000000000015500000000000000fb3378d51c",
    x"030b0000000000000155fffffffffffff50003e6831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f414c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2af31c",
    x"070a0000000000000155fffffffffffff8ef35fd731c",
    x"08020000000000000155fffffffffffff6f669e5d21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d78c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8571c",
    x"0209000000000000015500000000000000fb3378d01c",
    x"030b0000000000000155fffffffffffff50003e6841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2aec1c",
    x"070a0000000000000155fffffffffffff8ef35fd6f1c",
    x"08020000000000000155fffffffffffff6f669e5d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8581c",
    x"0209000000000000015500000000000000fb3378ca1c",
    x"030b0000000000000155fffffffffffff50003e6851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ae61c",
    x"070a0000000000000155fffffffffffff8ef35fd6c1c",
    x"08020000000000000155fffffffffffff6f669e5ce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe85a1c",
    x"0209000000000000015500000000000000fb3378c51c",
    x"030b0000000000000155fffffffffffff50003e6861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ae01c",
    x"070a0000000000000155fffffffffffff8ef35fd681c",
    x"08020000000000000155fffffffffffff6f669e5cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe85b1c",
    x"0209000000000000015500000000000000fb3378bf1c",
    x"030b0000000000000155fffffffffffff50003e6871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc0f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f413d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ada1c",
    x"070a0000000000000155fffffffffffff8ef35fd641c",
    x"08020000000000000155fffffffffffff6f669e5c91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d77b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe85c1c",
    x"0209000000000000015500000000000000fb3378b91c",
    x"030b0000000000000155fffffffffffff50003e6881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc0d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f413a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ad41c",
    x"070a0000000000000155fffffffffffff8ef35fd611c",
    x"08020000000000000155fffffffffffff6f669e5c61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe85d1c",
    x"0209000000000000015500000000000000fb3378b41c",
    x"030b0000000000000155fffffffffffff50003e6891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc0b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ace1c",
    x"070a0000000000000155fffffffffffff8ef35fd5d1c",
    x"08020000000000000155fffffffffffff6f669e5c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe85e1c",
    x"0209000000000000015500000000000000fb3378ae1c",
    x"030b0000000000000155fffffffffffff50003e68a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ac71c",
    x"070a0000000000000155fffffffffffff8ef35fd591c",
    x"08020000000000000155fffffffffffff6f669e5c21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d76f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe85f1c",
    x"0209000000000000015500000000000000fb3378a91c",
    x"030b0000000000000155fffffffffffff50003e68b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc061c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f412f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ac11c",
    x"070a0000000000000155fffffffffffff8ef35fd561c",
    x"08020000000000000155fffffffffffff6f669e5bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d76b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8601c",
    x"0209000000000000015500000000000000fb3378a31c",
    x"030b0000000000000155fffffffffffff50003e68c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f412b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2abb1c",
    x"070a0000000000000155fffffffffffff8ef35fd521c",
    x"08020000000000000155fffffffffffff6f669e5bd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8611c",
    x"0209000000000000015500000000000000fb33789d1c",
    x"030b0000000000000155fffffffffffff50003e68d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcc011c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2ab51c",
    x"070a0000000000000155fffffffffffff8ef35fd4f1c",
    x"08020000000000000155fffffffffffff6f669e5bb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8621c",
    x"0209000000000000015500000000000000fb3378981c",
    x"030b0000000000000155fffffffffffff50003e68e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcbfe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2aaf1c",
    x"070a0000000000000155fffffffffffff8ef35fd4b1c",
    x"08020000000000000155fffffffffffff6f669e5b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d75e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8641c",
    x"0209000000000000015500000000000000fb3378921c",
    x"030b0000000000000155fffffffffffff50003e68f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcbfc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2aa91c",
    x"070a0000000000000155fffffffffffff8ef35fd471c",
    x"08020000000000000155fffffffffffff6f669e5b61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d75a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8651c",
    x"0209000000000000015500000000000000fb33788d1c",
    x"030b0000000000000155fffffffffffff50003e6901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcbfa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f411c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2aa31c",
    x"070a0000000000000155fffffffffffff8ef35fd441c",
    x"08020000000000000155fffffffffffff6f669e5b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d7561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8661c",
    x"0209000000000000015500000000000000fb3378871c",
    x"030b0000000000000155fffffffffffff50003e6911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcbf71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f41181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd2a9c1c",
    x"070a0000000000000155fffffffffffff8ef35fd401c",
    x"08020000000000000155fffffffffffff6f669e5b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d7521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8671c",
    x"0209000000000000031f00000000000000fb3378811c",
    x"030b000000000000031ffffffffffffff50003e6921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcbf51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f41151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2a961c",
    x"070a000000000000031ffffffffffffff8ef35fd3d1c",
    x"0802000000000000031ffffffffffffff6f669e5af1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d74d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8681c",
    x"020900000000000000ae00000000000000fb33787c1c",
    x"030b00000000000000aefffffffffffff50003e6931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcbf21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f41111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2a901c",
    x"070a00000000000000aefffffffffffff8ef35fd391c",
    x"080200000000000000aefffffffffffff6f669e5ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d7491c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8691c",
    x"020900000000000001a400000000000000fb3378761c",
    x"030b00000000000001a4fffffffffffff50003e6941c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcbf01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f410d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2a8a1c",
    x"070a00000000000001a4fffffffffffff8ef35fd351c",
    x"080200000000000001a4fffffffffffff6f669e5aa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266d7451c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe86a1c",
    x"0209000000000000015600000000000000fb3378711c",
    x"030b0000000000000156fffffffffffff50003e6951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dcbee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f410a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd2a841c",
    x"070a0000000000000156fffffffffffff8ef35fd321c",
    x"08020000000000000156fffffffffffff6f669e5a71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d7411c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe86b1c",
    x"0209000000000000029500000000000000fb33786b1c",
    x"030b0000000000000295fffffffffffff50003e6961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcbeb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f41061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd2a7e1c",
    x"070a0000000000000295fffffffffffff8ef35fd2e1c",
    x"08020000000000000295fffffffffffff6f669e5a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d73d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe86c1c",
    x"0209000000000000029a00000000000000fb3378651c",
    x"030b000000000000029afffffffffffff50003e6971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcbe91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f41021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd2a781c",
    x"070a000000000000029afffffffffffff8ef35fd2a1c",
    x"0802000000000000029afffffffffffff6f669e5a31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe86d1c",
    x"020900000000000002aa00000000000000fb3378601c",
    x"030b00000000000002aafffffffffffff50003e6981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbe61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a711c",
    x"070a00000000000002aafffffffffffff8ef35fd271c",
    x"080200000000000002aafffffffffffff6f669e5a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe86f1c",
    x"020900000000000002aa00000000000000fb33785a1c",
    x"030b00000000000002aafffffffffffff50003e6991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbe41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a6b1c",
    x"070a00000000000002aafffffffffffff8ef35fd231c",
    x"080200000000000002aafffffffffffff6f669e59e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8701c",
    x"020900000000000002aa00000000000000fb3378551c",
    x"030b00000000000002aafffffffffffff50003e69a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbe21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40f71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a651c",
    x"070a00000000000002aafffffffffffff8ef35fd201c",
    x"080200000000000002aafffffffffffff6f669e59b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d72c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8711c",
    x"020900000000000002aa00000000000000fb33784f1c",
    x"030b00000000000002aafffffffffffff50003e69b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbdf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a5f1c",
    x"070a00000000000002aafffffffffffff8ef35fd1c1c",
    x"080200000000000002aafffffffffffff6f669e5991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8721c",
    x"020900000000000002aa00000000000000fb3378491c",
    x"030b00000000000002aafffffffffffff50003e69c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbdd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a591c",
    x"070a00000000000002aafffffffffffff8ef35fd181c",
    x"080200000000000002aafffffffffffff6f669e5971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8731c",
    x"020900000000000002aa00000000000000fb3378441c",
    x"030b00000000000002aafffffffffffff50003e69d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbda1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40ec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a531c",
    x"070a00000000000002aafffffffffffff8ef35fd151c",
    x"080200000000000002aafffffffffffff6f669e5941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d71f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8741c",
    x"020900000000000002aa00000000000000fb33783e1c",
    x"030b00000000000002aafffffffffffff50003e69e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbd81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a4c1c",
    x"070a00000000000002aafffffffffffff8ef35fd111c",
    x"080200000000000002aafffffffffffff6f669e5921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d71b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8751c",
    x"020900000000000002aa00000000000000fb3378391c",
    x"030b00000000000002aafffffffffffff50003e69f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbd51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40e51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a461c",
    x"070a00000000000002aafffffffffffff8ef35fd0d1c",
    x"080200000000000002aafffffffffffff6f669e5901c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8761c",
    x"020900000000000002aa00000000000000fb3378331c",
    x"030b00000000000002aafffffffffffff50003e6a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbd31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40e11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a401c",
    x"070a00000000000002aafffffffffffff8ef35fd0a1c",
    x"080200000000000002aafffffffffffff6f669e58d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7131c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8771c",
    x"020900000000000002aa00000000000000fb33782d1c",
    x"030b00000000000002aafffffffffffff50003e6a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbd11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a3a1c",
    x"070a00000000000002aafffffffffffff8ef35fd061c",
    x"080200000000000002aafffffffffffff6f669e58b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d70f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8791c",
    x"020900000000000002aa00000000000000fb3378281c",
    x"030b00000000000002aafffffffffffff50003e6a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40da1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a341c",
    x"070a00000000000002aafffffffffffff8ef35fd031c",
    x"080200000000000002aafffffffffffff6f669e5881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d70a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe87a1c",
    x"020900000000000002aa00000000000000fb3378221c",
    x"030b00000000000002aafffffffffffff50003e6a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbcc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40d61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a2e1c",
    x"070a00000000000002aafffffffffffff8ef35fcff1c",
    x"080200000000000002aafffffffffffff6f669e5861c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe87b1c",
    x"020900000000000002aa00000000000000fb33781d1c",
    x"030b00000000000002aafffffffffffff50003e6a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbc91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40d31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a281c",
    x"070a00000000000002aafffffffffffff8ef35fcfb1c",
    x"080200000000000002aafffffffffffff6f669e5841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d7021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe87c1c",
    x"020900000000000002aa00000000000000fb3378171c",
    x"030b00000000000002aafffffffffffff50003e6a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbc71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40cf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a211c",
    x"070a00000000000002aafffffffffffff8ef35fcf81c",
    x"080200000000000002aafffffffffffff6f669e5811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d6fe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe87d1c",
    x"0209000000000000031f00000000000000fb3378111c",
    x"030b000000000000031ffffffffffffff50003e6a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcbc51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f40cb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd2a1b1c",
    x"070a000000000000031ffffffffffffff8ef35fcf41c",
    x"0802000000000000031ffffffffffffff6f669e57f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d6fa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe87e1c",
    x"020900000000000000ae00000000000000fb33780c1c",
    x"030b00000000000000aefffffffffffff50003e6a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcbc21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f40c71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd2a151c",
    x"070a00000000000000aefffffffffffff8ef35fcf11c",
    x"080200000000000000aefffffffffffff6f669e57c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d6f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe87f1c",
    x"020900000000000001a400000000000000fb3378061c",
    x"030b00000000000001a4fffffffffffff50003e6a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcbc01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f40c41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd2a0f1c",
    x"070a00000000000001a4fffffffffffff8ef35fced1c",
    x"080200000000000001a4fffffffffffff6f669e57a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d6f11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe8801c",
    x"0209000000000000025600000000000000fb3378011c",
    x"030b0000000000000256fffffffffffff50003e6a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dcbbd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f40c01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd2a091c",
    x"070a0000000000000256fffffffffffff8ef35fce91c",
    x"08020000000000000256fffffffffffff6f669e5781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6ed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8811c",
    x"020900000000000002aa00000000000000fb3377fb1c",
    x"030b00000000000002aafffffffffffff50003e6aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbbb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40bc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd2a031c",
    x"070a00000000000002aafffffffffffff8ef35fce61c",
    x"080200000000000002aafffffffffffff6f669e5751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6e91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8831c",
    x"020900000000000002aa00000000000000fb3377f51c",
    x"030b00000000000002aafffffffffffff50003e6ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbb81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40b91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29fc1c",
    x"070a00000000000002aafffffffffffff8ef35fce21c",
    x"080200000000000002aafffffffffffff6f669e5731c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6e51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8841c",
    x"020900000000000002aa00000000000000fb3377f01c",
    x"030b00000000000002aafffffffffffff50003e6ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbb61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40b51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29f61c",
    x"070a00000000000002aafffffffffffff8ef35fcde1c",
    x"080200000000000002aafffffffffffff6f669e5701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8851c",
    x"020900000000000002aa00000000000000fb3377ea1c",
    x"030b00000000000002aafffffffffffff50003e6ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbb41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40b11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29f01c",
    x"070a00000000000002aafffffffffffff8ef35fcdb1c",
    x"080200000000000002aafffffffffffff6f669e56e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6dc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8861c",
    x"020900000000000002aa00000000000000fb3377e51c",
    x"030b00000000000002aafffffffffffff50003e6ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbb11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40ae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29ea1c",
    x"070a00000000000002aafffffffffffff8ef35fcd71c",
    x"080200000000000002aafffffffffffff6f669e56c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8871c",
    x"020900000000000002aa00000000000000fb3377df1c",
    x"030b00000000000002aafffffffffffff50003e6af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbaf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40aa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29e41c",
    x"070a00000000000002aafffffffffffff8ef35fcd41c",
    x"080200000000000002aafffffffffffff6f669e5691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6d41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8881c",
    x"020900000000000002aa00000000000000fb3377d91c",
    x"030b00000000000002aafffffffffffff50003e6b01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40a61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29de1c",
    x"070a00000000000002aafffffffffffff8ef35fcd01c",
    x"080200000000000002aafffffffffffff6f669e5671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6d01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8891c",
    x"020900000000000002aa00000000000000fb3377d41c",
    x"030b00000000000002aafffffffffffff50003e6b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcbaa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40a31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29d81c",
    x"070a00000000000002aafffffffffffff8ef35fccc1c",
    x"080200000000000002aafffffffffffff6f669e5651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6cc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe88a1c",
    x"020900000000000002aa00000000000000fb3377ce1c",
    x"030b00000000000002aafffffffffffff50003e6b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcba81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f409f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29d11c",
    x"070a00000000000002aafffffffffffff8ef35fcc91c",
    x"080200000000000002aafffffffffffff6f669e5621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe88b1c",
    x"020900000000000002aa00000000000000fb3377c91c",
    x"030b00000000000002aafffffffffffff50003e6b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcba51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f409b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29cb1c",
    x"070a00000000000002aafffffffffffff8ef35fcc51c",
    x"080200000000000002aafffffffffffff6f669e5601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe88c1c",
    x"020900000000000002aa00000000000000fb3377c31c",
    x"030b00000000000002aafffffffffffff50003e6b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcba31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29c51c",
    x"070a00000000000002aafffffffffffff8ef35fcc11c",
    x"080200000000000002aafffffffffffff6f669e55d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6bf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe88e1c",
    x"020900000000000002aa00000000000000fb3377bd1c",
    x"030b00000000000002aafffffffffffff50003e6b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcba01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29bf1c",
    x"070a00000000000002aafffffffffffff8ef35fcbe1c",
    x"080200000000000002aafffffffffffff6f669e55b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6bb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe88f1c",
    x"020900000000000002aa00000000000000fb3377b81c",
    x"030b00000000000002aafffffffffffff50003e6b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb9e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40901c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29b91c",
    x"070a00000000000002aafffffffffffff8ef35fcba1c",
    x"080200000000000002aafffffffffffff6f669e5591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6b71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8901c",
    x"020900000000000002aa00000000000000fb3377b21c",
    x"030b00000000000002aafffffffffffff50003e6b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb9b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f408d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29b31c",
    x"070a00000000000002aafffffffffffff8ef35fcb71c",
    x"080200000000000002aafffffffffffff6f669e5561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d6b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe8911c",
    x"0209000000000000029a00000000000000fb3377ad1c",
    x"030b000000000000029afffffffffffff50003e6b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dcb991c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f40891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd29ad1c",
    x"070a000000000000029afffffffffffff8ef35fcb31c",
    x"0802000000000000029afffffffffffff6f669e5541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8921c",
    x"020900000000000002aa00000000000000fb3377a71c",
    x"030b00000000000002aafffffffffffff50003e6b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40851c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29a61c",
    x"070a00000000000002aafffffffffffff8ef35fcaf1c",
    x"080200000000000002aafffffffffffff6f669e5511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d6aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8931c",
    x"0209000000000000031f00000000000000fb3377a11c",
    x"030b000000000000031ffffffffffffff50003e6b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcb941c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f40821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd29a01c",
    x"070a000000000000031ffffffffffffff8ef35fcac1c",
    x"0802000000000000031ffffffffffffff6f669e54f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d6a61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8941c",
    x"020900000000000000ae00000000000000fb33779c1c",
    x"030b00000000000000aefffffffffffff50003e6ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcb921c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f407e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd299a1c",
    x"070a00000000000000aefffffffffffff8ef35fca81c",
    x"080200000000000000aefffffffffffff6f669e54d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d6a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8951c",
    x"020900000000000001a400000000000000fb3377961c",
    x"030b00000000000001a4fffffffffffff50003e6bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcb8f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f407a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd29941c",
    x"070a00000000000001a4fffffffffffff8ef35fca41c",
    x"080200000000000001a4fffffffffffff6f669e54a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266d69d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe8961c",
    x"0209000000000000029600000000000000fb3377911c",
    x"030b0000000000000296fffffffffffff50003e6bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dcb8d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f40761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd298e1c",
    x"070a0000000000000296fffffffffffff8ef35fca11c",
    x"08020000000000000296fffffffffffff6f669e5481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d6991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe8981c",
    x"0209000000000000016a00000000000000fb33778b1c",
    x"030b000000000000016afffffffffffff50003e6bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcb8b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f40731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd29881c",
    x"070a000000000000016afffffffffffff8ef35fc9d1c",
    x"0802000000000000016afffffffffffff6f669e5451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266d6951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe8991c",
    x"020900000000000002a900000000000000fb3377851c",
    x"030b00000000000002a9fffffffffffff50003e6be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a9fffffffffffff4099dcb881c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f406f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd29811c",
    x"070a00000000000002a9fffffffffffff8ef35fc9a1c",
    x"080200000000000002a9fffffffffffff6f669e5431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe89a1c",
    x"020900000000000002aa00000000000000fb3377801c",
    x"030b00000000000002aafffffffffffff50003e6bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f406b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd297b1c",
    x"070a00000000000002aafffffffffffff8ef35fc961c",
    x"080200000000000002aafffffffffffff6f669e5411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d68d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe89b1c",
    x"020900000000000002aa00000000000000fb33777a1c",
    x"030b00000000000002aafffffffffffff50003e6c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29751c",
    x"070a00000000000002aafffffffffffff8ef35fc921c",
    x"080200000000000002aafffffffffffff6f669e53e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6891c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe89c1c",
    x"020900000000000002aa00000000000000fb3377751c",
    x"030b00000000000002aafffffffffffff50003e6c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd296f1c",
    x"070a00000000000002aafffffffffffff8ef35fc8f1c",
    x"080200000000000002aafffffffffffff6f669e53c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe89d1c",
    x"020900000000000002aa00000000000000fb33776f1c",
    x"030b00000000000002aafffffffffffff50003e6c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb7e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40601c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29691c",
    x"070a00000000000002aafffffffffffff8ef35fc8b1c",
    x"080200000000000002aafffffffffffff6f669e53a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe89e1c",
    x"020900000000000002aa00000000000000fb3377691c",
    x"030b00000000000002aafffffffffffff50003e6c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb7c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f405d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29631c",
    x"070a00000000000002aafffffffffffff8ef35fc871c",
    x"080200000000000002aafffffffffffff6f669e5371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d67c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe89f1c",
    x"020900000000000002aa00000000000000fb3377641c",
    x"030b00000000000002aafffffffffffff50003e6c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb7a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd295d1c",
    x"070a00000000000002aafffffffffffff8ef35fc841c",
    x"080200000000000002aafffffffffffff6f669e5351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a01c",
    x"020900000000000002aa00000000000000fb33775e1c",
    x"030b00000000000002aafffffffffffff50003e6c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29561c",
    x"070a00000000000002aafffffffffffff8ef35fc801c",
    x"080200000000000002aafffffffffffff6f669e5321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6741c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a21c",
    x"020900000000000002aa00000000000000fb3377591c",
    x"030b00000000000002aafffffffffffff50003e6c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29501c",
    x"070a00000000000002aafffffffffffff8ef35fc7d1c",
    x"080200000000000002aafffffffffffff6f669e5301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d66f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a31c",
    x"020900000000000002aa00000000000000fb3377531c",
    x"030b00000000000002aafffffffffffff50003e6c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb721c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f404e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd294a1c",
    x"070a00000000000002aafffffffffffff8ef35fc791c",
    x"080200000000000002aafffffffffffff6f669e52e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d66b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a41c",
    x"020900000000000002aa00000000000000fb33774d1c",
    x"030b00000000000002aafffffffffffff50003e6c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f404a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29441c",
    x"070a00000000000002aafffffffffffff8ef35fc751c",
    x"080200000000000002aafffffffffffff6f669e52b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a51c",
    x"020900000000000002aa00000000000000fb3377481c",
    x"030b00000000000002aafffffffffffff50003e6c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb6d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd293e1c",
    x"070a00000000000002aafffffffffffff8ef35fc721c",
    x"080200000000000002aafffffffffffff6f669e5291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a61c",
    x"020900000000000002aa00000000000000fb3377421c",
    x"030b00000000000002aafffffffffffff50003e6ca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb6b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f40431c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd29381c",
    x"070a00000000000002aafffffffffffff8ef35fc6e1c",
    x"080200000000000002aafffffffffffff6f669e5261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266d65f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe8a71c",
    x"0209000000000000019a00000000000000fb33773d1c",
    x"030b000000000000019afffffffffffff50003e6cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dcb691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f403f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd29311c",
    x"070a000000000000019afffffffffffff8ef35fc6a1c",
    x"0802000000000000019afffffffffffff6f669e5241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d65a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8a81c",
    x"020900000000000002aa00000000000000fb3377371c",
    x"030b00000000000002aafffffffffffff50003e6cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f403c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd292b1c",
    x"070a00000000000002aafffffffffffff8ef35fc671c",
    x"080200000000000002aafffffffffffff6f669e5221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d6561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8a91c",
    x"0209000000000000031f00000000000000fb3377311c",
    x"030b000000000000031ffffffffffffff50003e6cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcb641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f40381c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd29251c",
    x"070a000000000000031ffffffffffffff8ef35fc631c",
    x"0802000000000000031ffffffffffffff6f669e51f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d6521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8aa1c",
    x"020900000000000000ae00000000000000fb33772c1c",
    x"030b00000000000000aefffffffffffff50003e6ce1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcb611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f40341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd291f1c",
    x"070a00000000000000aefffffffffffff8ef35fc601c",
    x"080200000000000000aefffffffffffff6f669e51d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d64e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8ac1c",
    x"020900000000000001a400000000000000fb3377261c",
    x"030b00000000000001a4fffffffffffff50003e6cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcb5f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f40311c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd29191c",
    x"070a00000000000001a4fffffffffffff8ef35fc5c1c",
    x"080200000000000001a4fffffffffffff6f669e51a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266d64a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe8ad1c",
    x"0209000000000000019600000000000000fb3377211c",
    x"030b0000000000000196fffffffffffff50003e6d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dcb5d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f402d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000196ffffffffffffff04cd29131c",
    x"070a0000000000000196fffffffffffff8ef35fc581c",
    x"08020000000000000196fffffffffffff6f669e5181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8ae1c",
    x"0209000000000000015500000000000000fb33771b1c",
    x"030b0000000000000155fffffffffffff50003e6d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb5a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd290d1c",
    x"070a0000000000000155fffffffffffff8ef35fc551c",
    x"08020000000000000155fffffffffffff6f669e5161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6411c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8af1c",
    x"0209000000000000015500000000000000fb3377151c",
    x"030b0000000000000155fffffffffffff50003e6d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40261c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd29061c",
    x"070a0000000000000155fffffffffffff8ef35fc511c",
    x"08020000000000000155fffffffffffff6f669e5131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d63d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b01c",
    x"0209000000000000015500000000000000fb3377101c",
    x"030b0000000000000155fffffffffffff50003e6d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40221c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd29001c",
    x"070a0000000000000155fffffffffffff8ef35fc4d1c",
    x"08020000000000000155fffffffffffff6f669e5111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b11c",
    x"0209000000000000015500000000000000fb33770a1c",
    x"030b0000000000000155fffffffffffff50003e6d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f401e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28fa1c",
    x"070a0000000000000155fffffffffffff8ef35fc4a1c",
    x"08020000000000000155fffffffffffff6f669e50e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b21c",
    x"0209000000000000015500000000000000fb3377051c",
    x"030b0000000000000155fffffffffffff50003e6d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f401b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28f41c",
    x"070a0000000000000155fffffffffffff8ef35fc461c",
    x"08020000000000000155fffffffffffff6f669e50c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b31c",
    x"0209000000000000015500000000000000fb3376ff1c",
    x"030b0000000000000155fffffffffffff50003e6d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb4e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28ee1c",
    x"070a0000000000000155fffffffffffff8ef35fc431c",
    x"08020000000000000155fffffffffffff6f669e50a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d62c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b41c",
    x"0209000000000000015500000000000000fb3376f91c",
    x"030b0000000000000155fffffffffffff50003e6d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb4c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40131c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28e81c",
    x"070a0000000000000155fffffffffffff8ef35fc3f1c",
    x"08020000000000000155fffffffffffff6f669e5071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b51c",
    x"0209000000000000015500000000000000fb3376f41c",
    x"030b0000000000000155fffffffffffff50003e6d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f400f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28e11c",
    x"070a0000000000000155fffffffffffff8ef35fc3b1c",
    x"08020000000000000155fffffffffffff6f669e5051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b71c",
    x"0209000000000000015500000000000000fb3376ee1c",
    x"030b0000000000000155fffffffffffff50003e6d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f400c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28db1c",
    x"070a0000000000000155fffffffffffff8ef35fc381c",
    x"08020000000000000155fffffffffffff6f669e5031c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b81c",
    x"0209000000000000015500000000000000fb3376e91c",
    x"030b0000000000000155fffffffffffff50003e6da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40081c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28d51c",
    x"070a0000000000000155fffffffffffff8ef35fc341c",
    x"08020000000000000155fffffffffffff6f669e5001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d61c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8b91c",
    x"0209000000000000015500000000000000fb3376e31c",
    x"030b0000000000000155fffffffffffff50003e6db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40041c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28cf1c",
    x"070a0000000000000155fffffffffffff8ef35fc301c",
    x"08020000000000000155fffffffffffff6f669e4fe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8ba1c",
    x"0209000000000000015500000000000000fb3376dd1c",
    x"030b0000000000000155fffffffffffff50003e6dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb3f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f40011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28c91c",
    x"070a0000000000000155fffffffffffff8ef35fc2d1c",
    x"08020000000000000155fffffffffffff6f669e4fb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d6131c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8bb1c",
    x"0209000000000000015500000000000000fb3376d81c",
    x"030b0000000000000155fffffffffffff50003e6dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb3d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ffd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28c31c",
    x"070a0000000000000155fffffffffffff8ef35fc291c",
    x"08020000000000000155fffffffffffff6f669e4f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d60f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8bc1c",
    x"0209000000000000015500000000000000fb3376d21c",
    x"030b0000000000000155fffffffffffff50003e6de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb3b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ff91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28bd1c",
    x"070a0000000000000155fffffffffffff8ef35fc261c",
    x"08020000000000000155fffffffffffff6f669e4f71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266d60b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbe8bd1c",
    x"020900000000000002a500000000000000fb3376cd1c",
    x"030b00000000000002a5fffffffffffff50003e6df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dcb381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f3ff61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd28b61c",
    x"070a00000000000002a5fffffffffffff8ef35fc221c",
    x"080200000000000002a5fffffffffffff6f669e4f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d6071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8be1c",
    x"020900000000000002aa00000000000000fb3376c71c",
    x"030b00000000000002aafffffffffffff50003e6e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ff21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd28b01c",
    x"070a00000000000002aafffffffffffff8ef35fc1e1c",
    x"080200000000000002aafffffffffffff6f669e4f21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d6031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8bf1c",
    x"0209000000000000031f00000000000000fb3376c11c",
    x"030b000000000000031ffffffffffffff50003e6e11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcb331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3fee1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd28aa1c",
    x"070a000000000000031ffffffffffffff8ef35fc1b1c",
    x"0802000000000000031ffffffffffffff6f669e4ef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d5fe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8c11c",
    x"020900000000000000ae00000000000000fb3376bc1c",
    x"030b00000000000000aefffffffffffff50003e6e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcb311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3feb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd28a41c",
    x"070a00000000000000aefffffffffffff8ef35fc171c",
    x"080200000000000000aefffffffffffff6f669e4ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d5fa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8c21c",
    x"020900000000000001a400000000000000fb3376b61c",
    x"030b00000000000001a4fffffffffffff50003e6e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcb2f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3fe71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd289e1c",
    x"070a00000000000001a4fffffffffffff8ef35fc131c",
    x"080200000000000001a4fffffffffffff6f669e4eb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d5f61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbe8c31c",
    x"020900000000000002a600000000000000fb3376b11c",
    x"030b00000000000002a6fffffffffffff50003e6e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dcb2c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3fe31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd28981c",
    x"070a00000000000002a6fffffffffffff8ef35fc101c",
    x"080200000000000002a6fffffffffffff6f669e4e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d5f21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe8c41c",
    x"0209000000000000016a00000000000000fb3376ab1c",
    x"030b000000000000016afffffffffffff50003e6e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dcb2a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3fe01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd28911c",
    x"070a000000000000016afffffffffffff8ef35fc0c1c",
    x"0802000000000000016afffffffffffff6f669e4e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d5ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe8c51c",
    x"0209000000000000016600000000000000fb3376a51c",
    x"030b0000000000000166fffffffffffff50003e6e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dcb271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f3fdc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd288b1c",
    x"070a0000000000000166fffffffffffff8ef35fc091c",
    x"08020000000000000166fffffffffffff6f669e4e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5e91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8c61c",
    x"0209000000000000015500000000000000fb3376a01c",
    x"030b0000000000000155fffffffffffff50003e6e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fd81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28851c",
    x"070a0000000000000155fffffffffffff8ef35fc051c",
    x"08020000000000000155fffffffffffff6f669e4e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5e51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8c71c",
    x"0209000000000000015500000000000000fb33769a1c",
    x"030b0000000000000155fffffffffffff50003e6e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fd51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd287f1c",
    x"070a0000000000000155fffffffffffff8ef35fc011c",
    x"08020000000000000155fffffffffffff6f669e4df1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5e11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8c81c",
    x"0209000000000000015500000000000000fb3376951c",
    x"030b0000000000000155fffffffffffff50003e6e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fd11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28791c",
    x"070a0000000000000155fffffffffffff8ef35fbfe1c",
    x"08020000000000000155fffffffffffff6f669e4dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5dd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8c91c",
    x"0209000000000000015500000000000000fb33768f1c",
    x"030b0000000000000155fffffffffffff50003e6ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb1e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fcd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28731c",
    x"070a0000000000000155fffffffffffff8ef35fbfa1c",
    x"08020000000000000155fffffffffffff6f669e4da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5d91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8cb1c",
    x"0209000000000000015500000000000000fb3376891c",
    x"030b0000000000000155fffffffffffff50003e6eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb1b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd286d1c",
    x"070a0000000000000155fffffffffffff8ef35fbf61c",
    x"08020000000000000155fffffffffffff6f669e4d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5d51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8cc1c",
    x"0209000000000000015500000000000000fb3376841c",
    x"030b0000000000000155fffffffffffff50003e6ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fc61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28661c",
    x"070a0000000000000155fffffffffffff8ef35fbf31c",
    x"08020000000000000155fffffffffffff6f669e4d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5d01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8cd1c",
    x"0209000000000000015500000000000000fb33767e1c",
    x"030b0000000000000155fffffffffffff50003e6ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fc21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28601c",
    x"070a0000000000000155fffffffffffff8ef35fbef1c",
    x"08020000000000000155fffffffffffff6f669e4d31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5cc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8ce1c",
    x"0209000000000000015500000000000000fb3376791c",
    x"030b0000000000000155fffffffffffff50003e6ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fbf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd285a1c",
    x"070a0000000000000155fffffffffffff8ef35fbec1c",
    x"08020000000000000155fffffffffffff6f669e4d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5c81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8cf1c",
    x"0209000000000000015500000000000000fb3376731c",
    x"030b0000000000000155fffffffffffff50003e6ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fbb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28541c",
    x"070a0000000000000155fffffffffffff8ef35fbe81c",
    x"08020000000000000155fffffffffffff6f669e4ce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5c41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8d01c",
    x"0209000000000000015500000000000000fb33766d1c",
    x"030b0000000000000155fffffffffffff50003e6ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb0f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fb71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd284e1c",
    x"070a0000000000000155fffffffffffff8ef35fbe41c",
    x"08020000000000000155fffffffffffff6f669e4cc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5c01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8d11c",
    x"0209000000000000015500000000000000fb3376681c",
    x"030b0000000000000155fffffffffffff50003e6f01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb0d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fb41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28481c",
    x"070a0000000000000155fffffffffffff8ef35fbe11c",
    x"08020000000000000155fffffffffffff6f669e4c91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5bb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8d21c",
    x"0209000000000000015500000000000000fb3376621c",
    x"030b0000000000000155fffffffffffff50003e6f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcb0a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3fb01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28411c",
    x"070a0000000000000155fffffffffffff8ef35fbdd1c",
    x"08020000000000000155fffffffffffff6f669e4c71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d5b71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe8d31c",
    x"0209000000000000029500000000000000fb33765d1c",
    x"030b0000000000000295fffffffffffff50003e6f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcb081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3fac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd283b1c",
    x"070a0000000000000295fffffffffffff8ef35fbd91c",
    x"08020000000000000295fffffffffffff6f669e4c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5b31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8d51c",
    x"020900000000000002aa00000000000000fb3376571c",
    x"030b00000000000002aafffffffffffff50003e6f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcb051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3fa91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd28351c",
    x"070a00000000000002aafffffffffffff8ef35fbd61c",
    x"080200000000000002aafffffffffffff6f669e4c21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d5af1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8d61c",
    x"0209000000000000031f00000000000000fb3376511c",
    x"030b000000000000031ffffffffffffff50003e6f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcb031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3fa51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd282f1c",
    x"070a000000000000031ffffffffffffff8ef35fbd21c",
    x"0802000000000000031ffffffffffffff6f669e4c01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d5ab1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8d71c",
    x"020900000000000000ae00000000000000fb33764c1c",
    x"030b00000000000000aefffffffffffff50003e6f51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcb001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3fa11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd28291c",
    x"070a00000000000000aefffffffffffff8ef35fbcf1c",
    x"080200000000000000aefffffffffffff6f669e4bd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d5a61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8d81c",
    x"020900000000000001a400000000000000fb3376461c",
    x"030b00000000000001a4fffffffffffff50003e6f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcafe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3f9e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd28231c",
    x"070a00000000000001a4fffffffffffff8ef35fbcb1c",
    x"080200000000000001a4fffffffffffff6f669e4bb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266d5a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe8d91c",
    x"020900000000000001a600000000000000fb3376411c",
    x"030b00000000000001a6fffffffffffff50003e6f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dcafc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f3f9a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd281d1c",
    x"070a00000000000001a6fffffffffffff8ef35fbc71c",
    x"080200000000000001a6fffffffffffff6f669e4b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d59e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8da1c",
    x"0209000000000000015500000000000000fb33763b1c",
    x"030b0000000000000155fffffffffffff50003e6f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaf91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28161c",
    x"070a0000000000000155fffffffffffff8ef35fbc41c",
    x"08020000000000000155fffffffffffff6f669e4b61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d59a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8db1c",
    x"0209000000000000015500000000000000fb3376351c",
    x"030b0000000000000155fffffffffffff50003e6f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaf71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28101c",
    x"070a0000000000000155fffffffffffff8ef35fbc01c",
    x"08020000000000000155fffffffffffff6f669e4b41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5961c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8dc1c",
    x"0209000000000000015500000000000000fb3376301c",
    x"030b0000000000000155fffffffffffff50003e6fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaf41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f8f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd280a1c",
    x"070a0000000000000155fffffffffffff8ef35fbbc1c",
    x"08020000000000000155fffffffffffff6f669e4b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5921c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8dd1c",
    x"0209000000000000015500000000000000fb33762a1c",
    x"030b0000000000000155fffffffffffff50003e6fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaf21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f8b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd28041c",
    x"070a0000000000000155fffffffffffff8ef35fbb91c",
    x"08020000000000000155fffffffffffff6f669e4af1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d58d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8df1c",
    x"0209000000000000015500000000000000fb3376241c",
    x"030b0000000000000155fffffffffffff50003e6fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27fe1c",
    x"070a0000000000000155fffffffffffff8ef35fbb51c",
    x"08020000000000000155fffffffffffff6f669e4ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5891c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e01c",
    x"0209000000000000015500000000000000fb33761f1c",
    x"030b0000000000000155fffffffffffff50003e6fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27f81c",
    x"070a0000000000000155fffffffffffff8ef35fbb11c",
    x"08020000000000000155fffffffffffff6f669e4aa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5851c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e11c",
    x"0209000000000000015500000000000000fb3376191c",
    x"030b0000000000000155fffffffffffff50003e6fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcaeb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27f11c",
    x"070a0000000000000155fffffffffffff8ef35fbae1c",
    x"08020000000000000155fffffffffffff6f669e4a81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5811c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e21c",
    x"0209000000000000015500000000000000fb3376141c",
    x"030b0000000000000155fffffffffffff50003e6ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcae81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f7c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27eb1c",
    x"070a0000000000000155fffffffffffff8ef35fbaa1c",
    x"08020000000000000155fffffffffffff6f669e4a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d57d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e31c",
    x"0209000000000000015500000000000000fb33760e1c",
    x"030b0000000000000155fffffffffffff50003e7001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcae61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27e51c",
    x"070a0000000000000155fffffffffffff8ef35fba71c",
    x"08020000000000000155fffffffffffff6f669e4a31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e41c",
    x"0209000000000000015500000000000000fb3376081c",
    x"030b0000000000000155fffffffffffff50003e7011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcae31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27df1c",
    x"070a0000000000000155fffffffffffff8ef35fba31c",
    x"08020000000000000155fffffffffffff6f669e4a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5741c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e51c",
    x"0209000000000000015500000000000000fb3376031c",
    x"030b0000000000000155fffffffffffff50003e7021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcae11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27d91c",
    x"070a0000000000000155fffffffffffff8ef35fb9f1c",
    x"08020000000000000155fffffffffffff6f669e49e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5701c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e61c",
    x"0209000000000000015500000000000000fb3375fd1c",
    x"030b0000000000000155fffffffffffff50003e7031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcadf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f6e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27d31c",
    x"070a0000000000000155fffffffffffff8ef35fb9c1c",
    x"08020000000000000155fffffffffffff6f669e49c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d56c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e71c",
    x"0209000000000000015500000000000000fb3375f81c",
    x"030b0000000000000155fffffffffffff50003e7041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcadc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f6a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27cd1c",
    x"070a0000000000000155fffffffffffff8ef35fb981c",
    x"08020000000000000155fffffffffffff6f669e4991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d5681c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8e91c",
    x"0209000000000000015500000000000000fb3375f21c",
    x"030b0000000000000155fffffffffffff50003e7051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcada1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd27c61c",
    x"070a0000000000000155fffffffffffff8ef35fb941c",
    x"08020000000000000155fffffffffffff6f669e4971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d5631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe8ea1c",
    x"0209000000000000029500000000000000fb3375ec1c",
    x"030b0000000000000295fffffffffffff50003e7061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcad71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3f631c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd27c01c",
    x"070a0000000000000295fffffffffffff8ef35fb911c",
    x"08020000000000000295fffffffffffff6f669e4941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d55f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8eb1c",
    x"020900000000000002aa00000000000000fb3375e71c",
    x"030b00000000000002aafffffffffffff50003e7071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcad51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f5f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27ba1c",
    x"070a00000000000002aafffffffffffff8ef35fb8d1c",
    x"080200000000000002aafffffffffffff6f669e4921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d55b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe8ec1c",
    x"0209000000000000031f00000000000000fb3375e11c",
    x"030b000000000000031ffffffffffffff50003e7081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcad21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3f5b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd27b41c",
    x"070a000000000000031ffffffffffffff8ef35fb8a1c",
    x"0802000000000000031ffffffffffffff6f669e4901c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d5571c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe8ed1c",
    x"020900000000000000ae00000000000000fb3375dc1c",
    x"030b00000000000000aefffffffffffff50003e7091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dcad01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3f581c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd27ae1c",
    x"070a00000000000000aefffffffffffff8ef35fb861c",
    x"080200000000000000aefffffffffffff6f669e48d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d5531c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe8ee1c",
    x"020900000000000001a400000000000000fb3375d61c",
    x"030b00000000000001a4fffffffffffff50003e70a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dcace1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3f541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd27a81c",
    x"070a00000000000001a4fffffffffffff8ef35fb821c",
    x"080200000000000001a4fffffffffffff6f669e48b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d54f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe8ef1c",
    x"0209000000000000016600000000000000fb3375d01c",
    x"030b0000000000000166fffffffffffff50003e70b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dcacb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f3f501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd27a11c",
    x"070a0000000000000166fffffffffffff8ef35fb7f1c",
    x"08020000000000000166fffffffffffff6f669e4891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d54a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe8f01c",
    x"0209000000000000015500000000000000fb3375cb1c",
    x"030b0000000000000155fffffffffffff50003e70c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dcac91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3f4d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd279b1c",
    x"070a0000000000000155fffffffffffff8ef35fb7b1c",
    x"08020000000000000155fffffffffffff6f669e4861c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d5461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe8f11c",
    x"0209000000000000029500000000000000fb3375c51c",
    x"030b0000000000000295fffffffffffff50003e70d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dcac61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3f491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd27951c",
    x"070a0000000000000295fffffffffffff8ef35fb771c",
    x"08020000000000000295fffffffffffff6f669e4841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f31c",
    x"020900000000000002aa00000000000000fb3375c01c",
    x"030b00000000000002aafffffffffffff50003e70e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcac41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd278f1c",
    x"070a00000000000002aafffffffffffff8ef35fb741c",
    x"080200000000000002aafffffffffffff6f669e4811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d53e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f41c",
    x"020900000000000002aa00000000000000fb3375ba1c",
    x"030b00000000000002aafffffffffffff50003e70f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcac11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27891c",
    x"070a00000000000002aafffffffffffff8ef35fb701c",
    x"080200000000000002aafffffffffffff6f669e47f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d53a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f51c",
    x"020900000000000002aa00000000000000fb3375b41c",
    x"030b00000000000002aafffffffffffff50003e7101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcabf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f3e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27831c",
    x"070a00000000000002aafffffffffffff8ef35fb6d1c",
    x"080200000000000002aafffffffffffff6f669e47d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f61c",
    x"020900000000000002aa00000000000000fb3375af1c",
    x"030b00000000000002aafffffffffffff50003e7111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcabd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f3a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd277d1c",
    x"070a00000000000002aafffffffffffff8ef35fb691c",
    x"080200000000000002aafffffffffffff6f669e47a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f71c",
    x"020900000000000002aa00000000000000fb3375a91c",
    x"030b00000000000002aafffffffffffff50003e7121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcaba1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27761c",
    x"070a00000000000002aafffffffffffff8ef35fb651c",
    x"080200000000000002aafffffffffffff6f669e4781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d52d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f81c",
    x"020900000000000002aa00000000000000fb3375a41c",
    x"030b00000000000002aafffffffffffff50003e7131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcab81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f331c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27701c",
    x"070a00000000000002aafffffffffffff8ef35fb621c",
    x"080200000000000002aafffffffffffff6f669e4751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5291c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8f91c",
    x"020900000000000002aa00000000000000fb33759e1c",
    x"030b00000000000002aafffffffffffff50003e7141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcab51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f2f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd276a1c",
    x"070a00000000000002aafffffffffffff8ef35fb5e1c",
    x"080200000000000002aafffffffffffff6f669e4731c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5251c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8fa1c",
    x"020900000000000002aa00000000000000fb3375981c",
    x"030b00000000000002aafffffffffffff50003e7151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcab31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f2c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27641c",
    x"070a00000000000002aafffffffffffff8ef35fb5a1c",
    x"080200000000000002aafffffffffffff6f669e4711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8fb1c",
    x"020900000000000002aa00000000000000fb3375931c",
    x"030b00000000000002aafffffffffffff50003e7161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcab01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd275e1c",
    x"070a00000000000002aafffffffffffff8ef35fb571c",
    x"080200000000000002aafffffffffffff6f669e46e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d51c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8fd1c",
    x"020900000000000002aa00000000000000fb33758d1c",
    x"030b00000000000002aafffffffffffff50003e7161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcaae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27581c",
    x"070a00000000000002aafffffffffffff8ef35fb531c",
    x"080200000000000002aafffffffffffff6f669e46c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8fe1c",
    x"020900000000000002aa00000000000000fb3375881c",
    x"030b00000000000002aafffffffffffff50003e7171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcaac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f211c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27511c",
    x"070a00000000000002aafffffffffffff8ef35fb4f1c",
    x"080200000000000002aafffffffffffff6f669e4691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d5141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe8ff1c",
    x"020900000000000002aa00000000000000fb3375821c",
    x"030b00000000000002aafffffffffffff50003e7181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcaa91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f1d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd274b1c",
    x"070a00000000000002aafffffffffffff8ef35fb4c1c",
    x"080200000000000002aafffffffffffff6f669e4671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266d5101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe9001c",
    x"0209000000000000019a00000000000000fb33757c1c",
    x"030b000000000000019afffffffffffff50003e7191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dcaa71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f3f191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd27451c",
    x"070a000000000000019afffffffffffff8ef35fb481c",
    x"0802000000000000019afffffffffffff6f669e4651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d50c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9011c",
    x"020900000000000002aa00000000000000fb3375771c",
    x"030b00000000000002aafffffffffffff50003e71a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dcaa41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f161c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd273f1c",
    x"070a00000000000002aafffffffffffff8ef35fb451c",
    x"080200000000000002aafffffffffffff6f669e4621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d5071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9021c",
    x"0209000000000000031f00000000000000fb3375711c",
    x"030b000000000000031ffffffffffffff50003e71b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dcaa21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3f121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd27391c",
    x"070a000000000000031ffffffffffffff8ef35fb411c",
    x"0802000000000000031ffffffffffffff6f669e4601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d5031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9031c",
    x"020900000000000000ae00000000000000fb33756c1c",
    x"030b00000000000000aefffffffffffff50003e71c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dca9f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3f0e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd27331c",
    x"070a00000000000000aefffffffffffff8ef35fb3d1c",
    x"080200000000000000aefffffffffffff6f669e45d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d4ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9041c",
    x"020900000000000001a400000000000000fb3375661c",
    x"030b00000000000001a4fffffffffffff50003e71d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dca9d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3f0b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd272d1c",
    x"070a00000000000001a4fffffffffffff8ef35fb3a1c",
    x"080200000000000001a4fffffffffffff6f669e45b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d4fb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe9051c",
    x"0209000000000000026600000000000000fb3375601c",
    x"030b0000000000000266fffffffffffff50003e71e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dca9b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f3f071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000266ffffffffffffff04cd27261c",
    x"070a0000000000000266fffffffffffff8ef35fb361c",
    x"08020000000000000266fffffffffffff6f669e4591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4f71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9071c",
    x"020900000000000002aa00000000000000fb33755b1c",
    x"030b00000000000002aafffffffffffff50003e71f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27201c",
    x"070a00000000000002aafffffffffffff8ef35fb321c",
    x"080200000000000002aafffffffffffff6f669e4561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4f31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9081c",
    x"020900000000000002aa00000000000000fb3375551c",
    x"030b00000000000002aafffffffffffff50003e7201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3f001c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd271a1c",
    x"070a00000000000002aafffffffffffff8ef35fb2f1c",
    x"080200000000000002aafffffffffffff6f669e4541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9091c",
    x"020900000000000002aa00000000000000fb3375501c",
    x"030b00000000000002aafffffffffffff50003e7211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3efc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27141c",
    x"070a00000000000002aafffffffffffff8ef35fb2b1c",
    x"080200000000000002aafffffffffffff6f669e4511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4ea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe90a1c",
    x"020900000000000002aa00000000000000fb33754a1c",
    x"030b00000000000002aafffffffffffff50003e7221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ef81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd270e1c",
    x"070a00000000000002aafffffffffffff8ef35fb271c",
    x"080200000000000002aafffffffffffff6f669e44f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4e61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe90b1c",
    x"020900000000000002aa00000000000000fb3375441c",
    x"030b00000000000002aafffffffffffff50003e7231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca8e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ef51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27081c",
    x"070a00000000000002aafffffffffffff8ef35fb241c",
    x"080200000000000002aafffffffffffff6f669e44d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4e21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe90c1c",
    x"020900000000000002aa00000000000000fb33753f1c",
    x"030b00000000000002aafffffffffffff50003e7241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca8c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ef11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd27011c",
    x"070a00000000000002aafffffffffffff8ef35fb201c",
    x"080200000000000002aafffffffffffff6f669e44a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4de1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe90d1c",
    x"020900000000000002aa00000000000000fb3375391c",
    x"030b00000000000002aafffffffffffff50003e7251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca8a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3eed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26fb1c",
    x"070a00000000000002aafffffffffffff8ef35fb1d1c",
    x"080200000000000002aafffffffffffff6f669e4481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4d91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe90e1c",
    x"020900000000000002aa00000000000000fb3375341c",
    x"030b00000000000002aafffffffffffff50003e7261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3eea1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26f51c",
    x"070a00000000000002aafffffffffffff8ef35fb191c",
    x"080200000000000002aafffffffffffff6f669e4461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4d51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe90f1c",
    x"020900000000000002aa00000000000000fb33752e1c",
    x"030b00000000000002aafffffffffffff50003e7271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ee61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26ef1c",
    x"070a00000000000002aafffffffffffff8ef35fb151c",
    x"080200000000000002aafffffffffffff6f669e4431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4d11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9111c",
    x"020900000000000002aa00000000000000fb3375281c",
    x"030b00000000000002aafffffffffffff50003e7281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ee21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26e91c",
    x"070a00000000000002aafffffffffffff8ef35fb121c",
    x"080200000000000002aafffffffffffff6f669e4411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4cd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9121c",
    x"020900000000000002aa00000000000000fb3375231c",
    x"030b00000000000002aafffffffffffff50003e7291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3edf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26e31c",
    x"070a00000000000002aafffffffffffff8ef35fb0e1c",
    x"080200000000000002aafffffffffffff6f669e43e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4c91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9131c",
    x"020900000000000002aa00000000000000fb33751d1c",
    x"030b00000000000002aafffffffffffff50003e72a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca7d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3edb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26dc1c",
    x"070a00000000000002aafffffffffffff8ef35fb0a1c",
    x"080200000000000002aafffffffffffff6f669e43c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4c41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9141c",
    x"020900000000000002aa00000000000000fb3375181c",
    x"030b00000000000002aafffffffffffff50003e72b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca7b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ed71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26d61c",
    x"070a00000000000002aafffffffffffff8ef35fb071c",
    x"080200000000000002aafffffffffffff6f669e43a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4c01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9151c",
    x"020900000000000002aa00000000000000fb3375121c",
    x"030b00000000000002aafffffffffffff50003e72c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ed41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26d01c",
    x"070a00000000000002aafffffffffffff8ef35fb031c",
    x"080200000000000002aafffffffffffff6f669e4371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4bc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9161c",
    x"020900000000000002aa00000000000000fb33750c1c",
    x"030b00000000000002aafffffffffffff50003e72d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ed01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26ca1c",
    x"070a00000000000002aafffffffffffff8ef35fb001c",
    x"080200000000000002aafffffffffffff6f669e4351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4b81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9171c",
    x"020900000000000002aa00000000000000fb3375071c",
    x"030b00000000000002aafffffffffffff50003e72e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca741c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ecc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd26c41c",
    x"070a00000000000002aafffffffffffff8ef35fafc1c",
    x"080200000000000002aafffffffffffff6f669e4321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d4b41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9181c",
    x"0209000000000000031f00000000000000fb3375011c",
    x"030b000000000000031ffffffffffffff50003e72f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dca711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3ec91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd26be1c",
    x"070a000000000000031ffffffffffffff8ef35faf81c",
    x"0802000000000000031ffffffffffffff6f669e4301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d4b01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9191c",
    x"020900000000000000ae00000000000000fb3374fc1c",
    x"030b00000000000000aefffffffffffff50003e7301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dca6f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3ec51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd26b81c",
    x"070a00000000000000aefffffffffffff8ef35faf51c",
    x"080200000000000000aefffffffffffff6f669e42e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d4ab1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe91b1c",
    x"020900000000000001a400000000000000fb3374f61c",
    x"030b00000000000001a4fffffffffffff50003e7311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dca6c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3ec11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd26b11c",
    x"070a00000000000001a4fffffffffffff8ef35faf11c",
    x"080200000000000001a4fffffffffffff6f669e42b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d4a71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbe91c1c",
    x"020900000000000001aa00000000000000fb3374f01c",
    x"030b00000000000001aafffffffffffff50003e7321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dca6a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f3ebe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd26ab1c",
    x"070a00000000000001aafffffffffffff8ef35faed1c",
    x"080200000000000001aafffffffffffff6f669e4291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d4a31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe91d1c",
    x"0209000000000000029500000000000000fb3374eb1c",
    x"030b0000000000000295fffffffffffff50003e7331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dca671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3eba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd26a51c",
    x"070a0000000000000295fffffffffffff8ef35faea1c",
    x"08020000000000000295fffffffffffff6f669e4261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266d49f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe91e1c",
    x"0209000000000000015a00000000000000fb3374e51c",
    x"030b000000000000015afffffffffffff50003e7341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dca651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3eb61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd269f1c",
    x"070a000000000000015afffffffffffff8ef35fae61c",
    x"0802000000000000015afffffffffffff6f669e4241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d49b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe91f1c",
    x"0209000000000000025500000000000000fb3374e01c",
    x"030b0000000000000255fffffffffffff50003e7351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dca631c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f3eb31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd26991c",
    x"070a0000000000000255fffffffffffff8ef35fae21c",
    x"08020000000000000255fffffffffffff6f669e4221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266d4961c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe9201c",
    x"020900000000000002a900000000000000fb3374da1c",
    x"030b0000000000000155fffffffffffff50003e7361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dca601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3eaf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd26931c",
    x"070a0000000000000155fffffffffffff8ef35fadf1c",
    x"080200000000000002a9fffffffffffff6f669e41f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d4921c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9211c",
    x"0209000000000000029a00000000000000fb3374d41c",
    x"030b0000000000000265fffffffffffff50003e7371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dca5e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f3eab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd268c1c",
    x"070a0000000000000255fffffffffffff8ef35fadb1c",
    x"080200000000000002a9fffffffffffff6f669e41d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d48e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe9221c",
    x"0209000000000000015a00000000000000fb3374cf1c",
    x"030b0000000000000265fffffffffffff50003e7381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dca5b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ea81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd26861c",
    x"070a000000000000029afffffffffffff8ef35fad81c",
    x"0802000000000000019afffffffffffff6f669e41a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266d48a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe9231c",
    x"0209000000000000019900000000000000fb3374c91c",
    x"030b0000000000000166fffffffffffff50003e7391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dca591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f3ea41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd26801c",
    x"070a00000000000001a9fffffffffffff8ef35fad41c",
    x"0802000000000000026afffffffffffff6f669e4181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d4861c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002690000000000000b0bfbe9251c",
    x"0209000000000000016600000000000000fb3374c41c",
    x"030b00000000000001a6fffffffffffff50003e73a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dca561c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f3ea01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd267a1c",
    x"070a0000000000000199fffffffffffff8ef35fad01c",
    x"0802000000000000025afffffffffffff6f669e4161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266d4821c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9261c",
    x"0209000000000000015500000000000000fb3374be1c",
    x"030b000000000000015afffffffffffff50003e73a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dca541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3e9d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd26741c",
    x"070a000000000000016afffffffffffff8ef35facd1c",
    x"0802000000000000025afffffffffffff6f669e4131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d47d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe9271c",
    x"0209000000000000015a00000000000000fb3374b81c",
    x"030b0000000000000295fffffffffffff50003e73b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f3e991c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd266e1c",
    x"070a00000000000001aafffffffffffff8ef35fac91c",
    x"08020000000000000296fffffffffffff6f669e4111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266d4791c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002990000000000000b0bfbe9281c",
    x"020900000000000001a900000000000000fb3374b31c",
    x"030b0000000000000299fffffffffffff50003e73c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dca4f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3e951c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aaffffffffffffff04cd26681c",
    x"070a0000000000000165fffffffffffff8ef35fac51c",
    x"0802000000000000016afffffffffffff6f669e40e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266d4751c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe9291c",
    x"020900000000000002aa00000000000000fb3374ad1c",
    x"030b0000000000000169fffffffffffff50003e73d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dca4d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd26611c",
    x"070a00000000000002a9fffffffffffff8ef35fac21c",
    x"08020000000000000199fffffffffffff6f669e40c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000299ffffffffffffff0266d4711c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe92a1c",
    x"0209000000000000029a00000000000000fb3374a81c",
    x"030b000000000000019afffffffffffff50003e73e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dca4a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e8e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd265b1c",
    x"070a000000000000016afffffffffffff8ef35fabe1c",
    x"08020000000000000165fffffffffffff6f669e40a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266d46d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe92b1c",
    x"020900000000000002a600000000000000fb3374a21c",
    x"030b000000000000015afffffffffffff50003e73f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dca481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e8a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd26551c",
    x"070a000000000000025afffffffffffff8ef35faba1c",
    x"0802000000000000025afffffffffffff6f669e4071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266d4681c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe92c1c",
    x"020900000000000002aa00000000000000fb33749c1c",
    x"030b0000000000000265fffffffffffff50003e7401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dca451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001690000000000000b072f3e861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd264f1c",
    x"070a0000000000000159fffffffffffff8ef35fab71c",
    x"080200000000000001a9fffffffffffff6f669e4051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d4641c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe92d1c",
    x"0209000000000000015900000000000000fb3374971c",
    x"030b00000000000002a6fffffffffffff50003e7411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dca431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3e831c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd26491c",
    x"070a00000000000002a6fffffffffffff8ef35fab31c",
    x"0802000000000000016afffffffffffff6f669e4021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d4601c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe92f1c",
    x"0209000000000000031f00000000000000fb3374911c",
    x"030b000000000000031ffffffffffffff50003e7421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dca411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3e7f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd26431c",
    x"070a000000000000031ffffffffffffff8ef35fab01c",
    x"0802000000000000031ffffffffffffff6f669e4001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d45c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9301c",
    x"020900000000000000ae00000000000000fb33748c1c",
    x"030b00000000000000aefffffffffffff50003e7431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dca3e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3e7b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd263c1c",
    x"070a00000000000000aefffffffffffff8ef35faac1c",
    x"080200000000000000aefffffffffffff6f669e3fe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d4581c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9311c",
    x"020900000000000001a400000000000000fb3374861c",
    x"030b00000000000001a4fffffffffffff50003e7441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dca3c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3e781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd26361c",
    x"070a00000000000001a4fffffffffffff8ef35faa81c",
    x"080200000000000001a4fffffffffffff6f669e3fb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d4541c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe9321c",
    x"0209000000000000016a00000000000000fb3374801c",
    x"030b000000000000016afffffffffffff50003e7451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dca391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3e741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016affffffffffffff04cd26301c",
    x"070a000000000000016afffffffffffff8ef35faa51c",
    x"0802000000000000016afffffffffffff6f669e3f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d44f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9331c",
    x"0209000000000000015500000000000000fb33747b1c",
    x"030b0000000000000155fffffffffffff50003e7461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dca371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3e701c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd262a1c",
    x"070a0000000000000155fffffffffffff8ef35faa11c",
    x"08020000000000000155fffffffffffff6f669e3f71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266d44b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe9341c",
    x"0209000000000000019500000000000000fb3374751c",
    x"030b0000000000000195fffffffffffff50003e7471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dca341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f3e6d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd26241c",
    x"070a0000000000000195fffffffffffff8ef35fa9d1c",
    x"080200000000000002a5fffffffffffff6f669e3f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4471c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9351c",
    x"020900000000000002aa00000000000000fb33746f1c",
    x"030b00000000000002aafffffffffffff50003e7481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dca321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3e691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd261e1c",
    x"070a00000000000002aafffffffffffff8ef35fa9a1c",
    x"08020000000000000155fffffffffffff6f669e3f21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d4431c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbe9361c",
    x"0209000000000000029600000000000000fb33746a1c",
    x"030b00000000000001aafffffffffffff50003e7491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dca301c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3e651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd26171c",
    x"070a0000000000000256fffffffffffff8ef35fa961c",
    x"08020000000000000155fffffffffffff6f669e3ef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266d43f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe9371c",
    x"0209000000000000026500000000000000fb3374641c",
    x"030b00000000000002a9fffffffffffff50003e74a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dca2d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3e621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd26111c",
    x"070a000000000000029afffffffffffff8ef35fa921c",
    x"08020000000000000159fffffffffffff6f669e3ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266d43a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbe9391c",
    x"0209000000000000029600000000000000fb33745f1c",
    x"030b000000000000016afffffffffffff50003e74b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dca2b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3e5e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd260b1c",
    x"070a0000000000000159fffffffffffff8ef35fa8f1c",
    x"0802000000000000015afffffffffffff6f669e3eb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d4361c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe93a1c",
    x"0209000000000000016900000000000000fb3374591c",
    x"030b0000000000000295fffffffffffff50003e74c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dca281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e5a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019affffffffffffff04cd26051c",
    x"070a0000000000000196fffffffffffff8ef35fa8b1c",
    x"08020000000000000299fffffffffffff6f669e3e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d4321c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe93b1c",
    x"020900000000000002a500000000000000fb3374531c",
    x"030b0000000000000156fffffffffffff50003e74d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dca261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3e571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a5ffffffffffffff04cd25ff1c",
    x"070a00000000000002a6fffffffffffff8ef35fa871c",
    x"080200000000000001a5fffffffffffff6f669e3e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266d42e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe93c1c",
    x"0209000000000000025500000000000000fb33744e1c",
    x"030b000000000000016afffffffffffff50003e74e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dca231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f3e531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd25f91c",
    x"070a0000000000000295fffffffffffff8ef35fa841c",
    x"0802000000000000026afffffffffffff6f669e3e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d42a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe93d1c",
    x"0209000000000000029a00000000000000fb3374481c",
    x"030b0000000000000269fffffffffffff50003e74f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dca211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3e4f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd25f31c",
    x"070a0000000000000196fffffffffffff8ef35fa801c",
    x"08020000000000000165fffffffffffff6f669e3e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d4261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe93e1c",
    x"020900000000000001a600000000000000fb3374431c",
    x"030b000000000000019afffffffffffff50003e7501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dca1e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f3e4c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a6ffffffffffffff04cd25ec1c",
    x"070a000000000000026afffffffffffff8ef35fa7d1c",
    x"0802000000000000019afffffffffffff6f669e3df1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266d4211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbe93f1c",
    x"0209000000000000025a00000000000000fb33743d1c",
    x"030b00000000000002a9fffffffffffff50003e7511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dca1c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f3e481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a5ffffffffffffff04cd25e61c",
    x"070a00000000000002a6fffffffffffff8ef35fa791c",
    x"08020000000000000295fffffffffffff6f669e3dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d41d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbe9401c",
    x"0209000000000000029600000000000000fb3374371c",
    x"030b000000000000025afffffffffffff50003e7521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dca1a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f3e441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000165ffffffffffffff04cd25e01c",
    x"070a000000000000019afffffffffffff8ef35fa751c",
    x"0802000000000000029afffffffffffff6f669e3da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266d4191c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe9411c",
    x"0209000000000000019900000000000000fb3374321c",
    x"030b0000000000000156fffffffffffff50003e7531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dca171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f3e411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd25da1c",
    x"070a0000000000000166fffffffffffff8ef35fa721c",
    x"080200000000000001a9fffffffffffff6f669e3d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d4151c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe9431c",
    x"0209000000000000015600000000000000fb33742c1c",
    x"030b0000000000000169fffffffffffff50003e7541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dca151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f3e3d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd25d41c",
    x"070a0000000000000159fffffffffffff8ef35fa6e1c",
    x"08020000000000000255fffffffffffff6f669e3d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266d4111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9441c",
    x"0209000000000000029a00000000000000fb3374271c",
    x"030b00000000000002a9fffffffffffff50003e7551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dca121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3e391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd25ce1c",
    x"070a0000000000000159fffffffffffff8ef35fa6a1c",
    x"08020000000000000299fffffffffffff6f669e3d31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d40c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9451c",
    x"0209000000000000031f00000000000000fb3374211c",
    x"030b000000000000031ffffffffffffff50003e7561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dca101c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3e361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd25c71c",
    x"070a000000000000031ffffffffffffff8ef35fa671c",
    x"0802000000000000031ffffffffffffff6f669e3d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d4081c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9461c",
    x"020900000000000000ae00000000000000fb33741b1c",
    x"030b00000000000000aefffffffffffff50003e7571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dca0d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3e321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd25c11c",
    x"070a00000000000000aefffffffffffff8ef35fa631c",
    x"080200000000000000aefffffffffffff6f669e3ce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d4041c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9471c",
    x"020900000000000001a400000000000000fb3374161c",
    x"030b00000000000001a4fffffffffffff50003e7581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dca0b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3e2e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd25bb1c",
    x"070a00000000000001a4fffffffffffff8ef35fa5f1c",
    x"080200000000000001a4fffffffffffff6f669e3cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266d4001c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe9481c",
    x"0209000000000000026a00000000000000fb3374101c",
    x"030b000000000000026afffffffffffff50003e7591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dca091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f3e2b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026affffffffffffff04cd25b51c",
    x"070a000000000000026afffffffffffff8ef35fa5c1c",
    x"0802000000000000026afffffffffffff6f669e3c91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d3fc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9491c",
    x"0209000000000000015500000000000000fb33740b1c",
    x"030b0000000000000155fffffffffffff50003e7591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dca061c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f3e271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd25af1c",
    x"070a00000000000002a9fffffffffffff8ef35fa581c",
    x"08020000000000000155fffffffffffff6f669e3c71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d3f71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe94a1c",
    x"0209000000000000015500000000000000fb3374051c",
    x"030b0000000000000155fffffffffffff50003e75a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dca041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3e231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd25a91c",
    x"070a00000000000001aafffffffffffff8ef35fa551c",
    x"08020000000000000155fffffffffffff6f669e3c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266d3f31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe94b1c",
    x"0209000000000000015600000000000000fb3373ff1c",
    x"030b0000000000000155fffffffffffff50003e75b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dca011c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3e201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd25a21c",
    x"070a00000000000002aafffffffffffff8ef35fa511c",
    x"08020000000000000155fffffffffffff6f669e3c21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d3ef1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe94d1c",
    x"0209000000000000025500000000000000fb3373fa1c",
    x"030b0000000000000195fffffffffffff50003e75c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9ff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f3e1c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a9ffffffffffffff04cd259c1c",
    x"070a000000000000026afffffffffffff8ef35fa4d1c",
    x"08020000000000000195fffffffffffff6f669e3bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d3eb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe94e1c",
    x"0209000000000000016500000000000000fb3373f41c",
    x"030b00000000000002a9fffffffffffff50003e75d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc9fc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3e181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000259ffffffffffffff04cd25961c",
    x"070a0000000000000256fffffffffffff8ef35fa4a1c",
    x"08020000000000000299fffffffffffff6f669e3bd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d3e71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe94f1c",
    x"0209000000000000019900000000000000fb3373ef1c",
    x"030b0000000000000195fffffffffffff50003e75e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc9fa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd25901c",
    x"070a0000000000000266fffffffffffff8ef35fa461c",
    x"080200000000000002a6fffffffffffff6f669e3bb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d3e31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe9501c",
    x"0209000000000000016500000000000000fb3373e91c",
    x"030b0000000000000166fffffffffffff50003e75f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc9f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f3e111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd258a1c",
    x"070a0000000000000156fffffffffffff8ef35fa421c",
    x"0802000000000000025afffffffffffff6f669e3b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d3de1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe9511c",
    x"0209000000000000019500000000000000fb3373e31c",
    x"030b0000000000000265fffffffffffff50003e7601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc9f51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e0d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a9ffffffffffffff04cd25841c",
    x"070a000000000000025afffffffffffff8ef35fa3f1c",
    x"0802000000000000016afffffffffffff6f669e3b61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d3da1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe9521c",
    x"0209000000000000026a00000000000000fb3373de1c",
    x"030b00000000000002aafffffffffffff50003e7611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9f31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3e0a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000255ffffffffffffff04cd257e1c",
    x"070a0000000000000195fffffffffffff8ef35fa3b1c",
    x"08020000000000000195fffffffffffff6f669e3b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266d3d61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe9531c",
    x"0209000000000000025600000000000000fb3373d81c",
    x"030b00000000000002a5fffffffffffff50003e7621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dc9f01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3e061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000296ffffffffffffff04cd25771c",
    x"070a00000000000002a5fffffffffffff8ef35fa371c",
    x"08020000000000000295fffffffffffff6f669e3b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d3d21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe9541c",
    x"020900000000000001a900000000000000fb3373d31c",
    x"030b0000000000000155fffffffffffff50003e7631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc9ee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f3e021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd25711c",
    x"070a0000000000000256fffffffffffff8ef35fa341c",
    x"08020000000000000199fffffffffffff6f669e3af1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d3ce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe9551c",
    x"0209000000000000029500000000000000fb3373cd1c",
    x"030b0000000000000299fffffffffffff50003e7641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3dff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd256b1c",
    x"070a0000000000000266fffffffffffff8ef35fa301c",
    x"08020000000000000166fffffffffffff6f669e3ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d3c91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbe9571c",
    x"0209000000000000016900000000000000fb3373c71c",
    x"030b000000000000016afffffffffffff50003e7651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc9e91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f3dfb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a6ffffffffffffff04cd25651c",
    x"070a0000000000000256fffffffffffff8ef35fa2c1c",
    x"08020000000000000199fffffffffffff6f669e3aa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266d3c51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe9581c",
    x"0209000000000000026a00000000000000fb3373c21c",
    x"030b000000000000016afffffffffffff50003e7661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc9e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3df71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000256ffffffffffffff04cd255f1c",
    x"070a00000000000001a5fffffffffffff8ef35fa291c",
    x"08020000000000000266fffffffffffff6f669e3a71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d3c11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe9591c",
    x"020900000000000001a900000000000000fb3373bc1c",
    x"030b000000000000026afffffffffffff50003e7671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc9e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f3df41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000166ffffffffffffff04cd25591c",
    x"070a0000000000000166fffffffffffff8ef35fa251c",
    x"08020000000000000296fffffffffffff6f669e3a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266d3bd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe95a1c",
    x"020900000000000002a600000000000000fb3373b71c",
    x"030b000000000000015afffffffffffff50003e7681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc9e21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3df01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000299ffffffffffffff04cd25521c",
    x"070a0000000000000295fffffffffffff8ef35fa221c",
    x"080200000000000002a5fffffffffffff6f669e3a31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d3b91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe95b1c",
    x"0209000000000000031f00000000000000fb3373b11c",
    x"030b000000000000031ffffffffffffff50003e7691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc9df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3dec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd254c1c",
    x"070a000000000000031ffffffffffffff8ef35fa1e1c",
    x"0802000000000000031ffffffffffffff6f669e3a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d3b51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe95c1c",
    x"020900000000000000ae00000000000000fb3373ab1c",
    x"030b00000000000000aefffffffffffff50003e76a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc9dd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3de91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd25461c",
    x"070a00000000000000aefffffffffffff8ef35fa1a1c",
    x"080200000000000000aefffffffffffff6f669e39e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d3b01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe95d1c",
    x"020900000000000001a400000000000000fb3373a61c",
    x"030b00000000000001a4fffffffffffff50003e76b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc9da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3de51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd25401c",
    x"070a00000000000001a4fffffffffffff8ef35fa171c",
    x"080200000000000001a4fffffffffffff6f669e39c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266d3ac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbe95e1c",
    x"0209000000000000015a00000000000000fb3373a01c",
    x"030b000000000000015afffffffffffff50003e76c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc9d81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3de11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd253a1c",
    x"070a000000000000015afffffffffffff8ef35fa131c",
    x"0802000000000000015afffffffffffff6f669e3991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3a81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9601c",
    x"020900000000000001aa00000000000000fb33739b1c",
    x"030b0000000000000255fffffffffffff50003e76d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9d51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3dde1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd25341c",
    x"070a0000000000000155fffffffffffff8ef35fa0f1c",
    x"08020000000000000155fffffffffffff6f669e3971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266d3a41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbe9611c",
    x"0209000000000000016900000000000000fb3373951c",
    x"030b0000000000000269fffffffffffff50003e76e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc9d31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3dda1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd252d1c",
    x"070a00000000000002a6fffffffffffff8ef35fa0c1c",
    x"080200000000000001a5fffffffffffff6f669e3941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266d3a01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbe9621c",
    x"020900000000000001a600000000000000fb33738f1c",
    x"030b0000000000000296fffffffffffff50003e76f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc9d11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f3dd61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd25271c",
    x"070a000000000000029afffffffffffff8ef35fa081c",
    x"08020000000000000196fffffffffffff6f669e3921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266d39b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe9631c",
    x"0209000000000000026900000000000000fb33738a1c",
    x"030b0000000000000255fffffffffffff50003e7701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc9ce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f3dd31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000199ffffffffffffff04cd25211c",
    x"070a0000000000000265fffffffffffff8ef35fa041c",
    x"08020000000000000256fffffffffffff6f669e3901c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3971c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe9641c",
    x"0209000000000000015600000000000000fb3373841c",
    x"030b0000000000000155fffffffffffff50003e7711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f3dcf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000156ffffffffffffff04cd251b1c",
    x"070a00000000000002aafffffffffffff8ef35fa011c",
    x"08020000000000000155fffffffffffff6f669e38d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9651c",
    x"0209000000000000015500000000000000fb33737f1c",
    x"030b0000000000000155fffffffffffff50003e7721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9c91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3dcb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd25151c",
    x"070a00000000000002aafffffffffffff8ef35f9fd1c",
    x"08020000000000000155fffffffffffff6f669e38b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d38f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9661c",
    x"0209000000000000015500000000000000fb3373791c",
    x"030b0000000000000155fffffffffffff50003e7731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3dc81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd250f1c",
    x"070a00000000000002aafffffffffffff8ef35f9fa1c",
    x"08020000000000000155fffffffffffff6f669e3881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d38b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9671c",
    x"0209000000000000015500000000000000fb3373731c",
    x"030b0000000000000155fffffffffffff50003e7741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9c41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3dc41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd25091c",
    x"070a00000000000002aafffffffffffff8ef35f9f61c",
    x"08020000000000000155fffffffffffff6f669e3861c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9681c",
    x"0209000000000000015500000000000000fb33736e1c",
    x"030b0000000000000155fffffffffffff50003e7751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3dc11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd25021c",
    x"070a00000000000002aafffffffffffff8ef35f9f21c",
    x"08020000000000000155fffffffffffff6f669e3841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266d3821c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbe96a1c",
    x"0209000000000000025900000000000000fb3373681c",
    x"030b0000000000000259fffffffffffff50003e7751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc9bf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f3dbd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000259ffffffffffffff04cd24fc1c",
    x"070a00000000000001a6fffffffffffff8ef35f9ef1c",
    x"08020000000000000259fffffffffffff6f669e3811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d37e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe96b1c",
    x"0209000000000000015500000000000000fb3373631c",
    x"030b0000000000000155fffffffffffff50003e7761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3db91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd24f61c",
    x"070a00000000000002aafffffffffffff8ef35f9eb1c",
    x"08020000000000000155fffffffffffff6f669e37f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d37a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe96c1c",
    x"0209000000000000015500000000000000fb33735d1c",
    x"030b0000000000000155fffffffffffff50003e7771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3db61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000155ffffffffffffff04cd24f01c",
    x"070a00000000000002aafffffffffffff8ef35f9e71c",
    x"08020000000000000155fffffffffffff6f669e37c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d3761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbe96d1c",
    x"0209000000000000015900000000000000fb3373571c",
    x"030b0000000000000159fffffffffffff50003e7781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc9b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3db21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000159ffffffffffffff04cd24ea1c",
    x"070a00000000000002a6fffffffffffff8ef35f9e41c",
    x"08020000000000000159fffffffffffff6f669e37a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266d3721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe96e1c",
    x"0209000000000000016a00000000000000fb3373521c",
    x"030b0000000000000155fffffffffffff50003e7791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc9b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f3dae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000295ffffffffffffff04cd24e41c",
    x"070a0000000000000265fffffffffffff8ef35f9e01c",
    x"0802000000000000015afffffffffffff6f669e3781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266d36d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbe96f1c",
    x"0209000000000000015500000000000000fb33734c1c",
    x"030b0000000000000155fffffffffffff50003e77a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f3dab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015affffffffffffff04cd24dd1c",
    x"070a000000000000025afffffffffffff8ef35f9dc1c",
    x"08020000000000000195fffffffffffff6f669e3751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d3691c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbe9701c",
    x"020900000000000002aa00000000000000fb3373461c",
    x"030b00000000000002aafffffffffffff50003e77b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc9b11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3da71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"06180000000000000169ffffffffffffff04cd24d71c",
    x"070a0000000000000155fffffffffffff8ef35f9d91c",
    x"080200000000000002aafffffffffffff6f669e3731c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d3651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9711c",
    x"0209000000000000031f00000000000000fb3373411c",
    x"030b000000000000031ffffffffffffff50003e77c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc9ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3da31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031fffffffffffffff04cd24d11c",
    x"070a000000000000031ffffffffffffff8ef35f9d51c",
    x"0802000000000000031ffffffffffffff6f669e3701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d3611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9721c",
    x"020900000000000000ae00000000000000fb33733b1c",
    x"030b00000000000000aefffffffffffff50003e77d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc9ac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3da01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000aeffffffffffffff04cd24cb1c",
    x"070a00000000000000aefffffffffffff8ef35f9d11c",
    x"080200000000000000aefffffffffffff6f669e36e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d35d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9741c",
    x"020900000000000001a400000000000000fb3373361c",
    x"030b00000000000001a4fffffffffffff50003e77e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc9aa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3d9c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a4ffffffffffffff04cd24c51c",
    x"070a00000000000001a4fffffffffffff8ef35f9ce1c",
    x"080200000000000001a4fffffffffffff6f669e36c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266d3591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbe9751c",
    x"0209000000000000025a00000000000000fb3373301c",
    x"030b000000000000025afffffffffffff50003e77f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc9a71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f3d981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025affffffffffffff04cd24bf1c",
    x"070a000000000000025afffffffffffff8ef35f9ca1c",
    x"0802000000000000025afffffffffffff6f669e3691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3541c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9761c",
    x"020900000000000002aa00000000000000fb33732a1c",
    x"030b00000000000002aafffffffffffff50003e7801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9a51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d951c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd24b81c",
    x"070a00000000000002aafffffffffffff8ef35f9c61c",
    x"080200000000000002aafffffffffffff6f669e3671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d3501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe9771c",
    x"0209000000000000029a00000000000000fb3373251c",
    x"030b000000000000029afffffffffffff50003e7811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc9a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f3d911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029affffffffffffff04cd24b21c",
    x"070a000000000000029afffffffffffff8ef35f9c31c",
    x"0802000000000000029afffffffffffff6f669e3641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d34c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9781c",
    x"020900000000000002aa00000000000000fb33731f1c",
    x"030b00000000000002aafffffffffffff50003e7821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9a01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d8d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd24ac1c",
    x"070a00000000000002aafffffffffffff8ef35f9bf1c",
    x"080200000000000002aafffffffffffff6f669e3621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9791c",
    x"020900000000000002aa00000000000000fb33731a1c",
    x"030b00000000000002aafffffffffffff50003e7831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc99d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d8a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd24a61c",
    x"070a00000000000002aafffffffffffff8ef35f9bc1c",
    x"080200000000000002aafffffffffffff6f669e3601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe97a1c",
    x"020900000000000002aa00000000000000fb3373141c",
    x"030b00000000000002aafffffffffffff50003e7841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc99b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd24a01c",
    x"070a00000000000002aafffffffffffff8ef35f9b81c",
    x"080200000000000002aafffffffffffff6f669e35d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d33f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe97b1c",
    x"020900000000000002aa00000000000000fb33730e1c",
    x"030b00000000000002aafffffffffffff50003e7851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd249a1c",
    x"070a00000000000002aafffffffffffff8ef35f9b41c",
    x"080200000000000002aafffffffffffff6f669e35b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d33b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe97c1c",
    x"020900000000000002aa00000000000000fb3373091c",
    x"030b00000000000002aafffffffffffff50003e7861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d7f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd24941c",
    x"070a00000000000002aafffffffffffff8ef35f9b11c",
    x"080200000000000002aafffffffffffff6f669e3581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe97e1c",
    x"020900000000000002aa00000000000000fb3373031c",
    x"030b00000000000002aafffffffffffff50003e7871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9941c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d7b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd248d1c",
    x"070a00000000000002aafffffffffffff8ef35f9ad1c",
    x"080200000000000002aafffffffffffff6f669e3561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d3331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe97f1c",
    x"020900000000000002aa00000000000000fb3372fe1c",
    x"030b00000000000002aafffffffffffff50003e7881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc9911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3d771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aaffffffffffffff04cd24871c",
    x"070a00000000000002aafffffffffffff8ef35f9a91c",
    x"080200000000000002aafffffffffffff6f669e3541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d32f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbe9801c",
    x"0209000000000000016600000000000000fb3372f81c",
    x"030b0000000000000166fffffffffffff50003e7891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc98f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f3d741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd24811c",
    x"070a0000000000000166fffffffffffff8ef35f9a61c",
    x"08020000000000000166fffffffffffff6f669e3511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d32b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9811c",
    x"0209000000000000015500000000000000fb3372f21c",
    x"030b0000000000000155fffffffffffff50003e78a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc98c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d701c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd247b1c",
    x"070a0000000000000155fffffffffffff8ef35f9a21c",
    x"08020000000000000155fffffffffffff6f669e34f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d3261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9821c",
    x"0209000000000000015500000000000000fb3372ed1c",
    x"030b0000000000000155fffffffffffff50003e78b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc98a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d6c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24751c",
    x"070a0000000000000155fffffffffffff8ef35f99e1c",
    x"08020000000000000155fffffffffffff6f669e34c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d3221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9831c",
    x"0209000000000000015500000000000000fb3372e71c",
    x"030b0000000000000155fffffffffffff50003e78c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd246f1c",
    x"070a0000000000000155fffffffffffff8ef35f99b1c",
    x"08020000000000000155fffffffffffff6f669e34a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d31e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9841c",
    x"0209000000000000015500000000000000fb3372e21c",
    x"030b0000000000000155fffffffffffff50003e78d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24681c",
    x"070a0000000000000155fffffffffffff8ef35f9971c",
    x"08020000000000000155fffffffffffff6f669e3481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d31a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9851c",
    x"0209000000000000015500000000000000fb3372dc1c",
    x"030b0000000000000155fffffffffffff50003e78e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24621c",
    x"070a0000000000000155fffffffffffff8ef35f9931c",
    x"08020000000000000155fffffffffffff6f669e3451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266d3161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbe9871c",
    x"0209000000000000015900000000000000fb3372d61c",
    x"030b0000000000000159fffffffffffff50003e78f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc9801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f3d5e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd245c1c",
    x"070a0000000000000159fffffffffffff8ef35f9901c",
    x"08020000000000000159fffffffffffff6f669e3431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d3111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9881c",
    x"0209000000000000031f00000000000000fb3372d11c",
    x"030b000000000000031ffffffffffffff50003e78f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc97e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3d5a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd24561c",
    x"070a000000000000031ffffffffffffff8ef35f98c1c",
    x"0802000000000000031ffffffffffffff6f669e3401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d30d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9891c",
    x"020900000000000000ae00000000000000fb3372cb1c",
    x"030b00000000000000aefffffffffffff50003e7901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc97b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3d561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd24501c",
    x"070a00000000000000aefffffffffffff8ef35f9891c",
    x"080200000000000000aefffffffffffff6f669e33e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d3091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe98a1c",
    x"020900000000000001a400000000000000fb3372c61c",
    x"030b00000000000001a4fffffffffffff50003e7911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc9791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3d531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd244a1c",
    x"070a00000000000001a4fffffffffffff8ef35f9851c",
    x"080200000000000001a4fffffffffffff6f669e33c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d3051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe98b1c",
    x"0209000000000000029a00000000000000fb3372c01c",
    x"030b000000000000029afffffffffffff50003e7921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc9761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f3d4f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd24431c",
    x"070a000000000000029afffffffffffff8ef35f9811c",
    x"0802000000000000029afffffffffffff6f669e3391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d3011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe98c1c",
    x"0209000000000000016a00000000000000fb3372ba1c",
    x"030b000000000000016afffffffffffff50003e7931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc9741c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3d4b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd243d1c",
    x"070a000000000000016afffffffffffff8ef35f97e1c",
    x"0802000000000000016afffffffffffff6f669e3371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266d2fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe98d1c",
    x"0209000000000000016500000000000000fb3372b51c",
    x"030b0000000000000165fffffffffffff50003e7941c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc9711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f3d481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd24371c",
    x"070a0000000000000165fffffffffffff8ef35f97a1c",
    x"08020000000000000165fffffffffffff6f669e3341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2f81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe98e1c",
    x"0209000000000000015500000000000000fb3372af1c",
    x"030b0000000000000155fffffffffffff50003e7951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc96f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24311c",
    x"070a0000000000000155fffffffffffff8ef35f9761c",
    x"08020000000000000155fffffffffffff6f669e3321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2f41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe98f1c",
    x"0209000000000000015500000000000000fb3372aa1c",
    x"030b0000000000000155fffffffffffff50003e7961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc96c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd242b1c",
    x"070a0000000000000155fffffffffffff8ef35f9731c",
    x"08020000000000000155fffffffffffff6f669e3301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2f01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9911c",
    x"0209000000000000015500000000000000fb3372a41c",
    x"030b0000000000000155fffffffffffff50003e7971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc96a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d3d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24251c",
    x"070a0000000000000155fffffffffffff8ef35f96f1c",
    x"08020000000000000155fffffffffffff6f669e32d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9921c",
    x"0209000000000000015500000000000000fb33729e1c",
    x"030b0000000000000155fffffffffffff50003e7981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9681c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd241e1c",
    x"070a0000000000000155fffffffffffff8ef35f96b1c",
    x"08020000000000000155fffffffffffff6f669e32b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9931c",
    x"0209000000000000015500000000000000fb3372991c",
    x"030b0000000000000155fffffffffffff50003e7991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24181c",
    x"070a0000000000000155fffffffffffff8ef35f9681c",
    x"08020000000000000155fffffffffffff6f669e3281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2e31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9941c",
    x"0209000000000000015500000000000000fb3372931c",
    x"030b0000000000000155fffffffffffff50003e79a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9631c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24121c",
    x"070a0000000000000155fffffffffffff8ef35f9641c",
    x"08020000000000000155fffffffffffff6f669e3261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2df1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9951c",
    x"0209000000000000015500000000000000fb33728e1c",
    x"030b0000000000000155fffffffffffff50003e79b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d2e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd240c1c",
    x"070a0000000000000155fffffffffffff8ef35f9601c",
    x"08020000000000000155fffffffffffff6f669e3241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2db1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9961c",
    x"0209000000000000015500000000000000fb3372881c",
    x"030b0000000000000155fffffffffffff50003e79c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc95e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d2a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24061c",
    x"070a0000000000000155fffffffffffff8ef35f95d1c",
    x"08020000000000000155fffffffffffff6f669e3211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2d71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9971c",
    x"0209000000000000015500000000000000fb3372821c",
    x"030b0000000000000155fffffffffffff50003e79d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc95b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd24001c",
    x"070a0000000000000155fffffffffffff8ef35f9591c",
    x"08020000000000000155fffffffffffff6f669e31f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9981c",
    x"0209000000000000015500000000000000fb33727d1c",
    x"030b0000000000000155fffffffffffff50003e79e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23fa1c",
    x"070a0000000000000155fffffffffffff8ef35f9551c",
    x"08020000000000000155fffffffffffff6f669e31c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9991c",
    x"0209000000000000015500000000000000fb3372771c",
    x"030b0000000000000155fffffffffffff50003e79f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d1f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23f31c",
    x"070a0000000000000155fffffffffffff8ef35f9521c",
    x"08020000000000000155fffffffffffff6f669e31a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2ca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe99b1c",
    x"0209000000000000015500000000000000fb3372721c",
    x"030b0000000000000155fffffffffffff50003e7a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d1c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23ed1c",
    x"070a0000000000000155fffffffffffff8ef35f94e1c",
    x"08020000000000000155fffffffffffff6f669e3181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266d2c61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbe99c1c",
    x"0209000000000000016500000000000000fb33726c1c",
    x"030b0000000000000165fffffffffffff50003e7a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc9521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f3d181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd23e71c",
    x"070a0000000000000165fffffffffffff8ef35f94b1c",
    x"08020000000000000165fffffffffffff6f669e3151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2c21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe99d1c",
    x"0209000000000000015500000000000000fb3372661c",
    x"030b0000000000000155fffffffffffff50003e7a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc94f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23e11c",
    x"070a0000000000000155fffffffffffff8ef35f9471c",
    x"08020000000000000155fffffffffffff6f669e3131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d2be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe99e1c",
    x"0209000000000000031f00000000000000fb3372611c",
    x"030b000000000000031ffffffffffffff50003e7a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc94d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3d111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd23db1c",
    x"070a000000000000031ffffffffffffff8ef35f9431c",
    x"0802000000000000031ffffffffffffff6f669e3111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d2ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe99f1c",
    x"020900000000000000ae00000000000000fb33725b1c",
    x"030b00000000000000aefffffffffffff50003e7a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc94a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3d0d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd23d51c",
    x"070a00000000000000aefffffffffffff8ef35f9401c",
    x"080200000000000000aefffffffffffff6f669e30e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d2b51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9a01c",
    x"020900000000000001a400000000000000fb3372551c",
    x"030b00000000000001a4fffffffffffff50003e7a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc9481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3d091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd23ce1c",
    x"070a00000000000001a4fffffffffffff8ef35f93c1c",
    x"080200000000000001a4fffffffffffff6f669e30c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266d2b11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbe9a11c",
    x"0209000000000000019a00000000000000fb3372501c",
    x"030b000000000000019afffffffffffff50003e7a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc9451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f3d061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd23c81c",
    x"070a000000000000019afffffffffffff8ef35f9381c",
    x"0802000000000000019afffffffffffff6f669e3091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2ad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a21c",
    x"0209000000000000015500000000000000fb33724a1c",
    x"030b0000000000000155fffffffffffff50003e7a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3d021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23c21c",
    x"070a0000000000000155fffffffffffff8ef35f9351c",
    x"08020000000000000155fffffffffffff6f669e3071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2a91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a41c",
    x"0209000000000000015500000000000000fb3372451c",
    x"030b0000000000000155fffffffffffff50003e7a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cfe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23bc1c",
    x"070a0000000000000155fffffffffffff8ef35f9311c",
    x"08020000000000000155fffffffffffff6f669e3051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a51c",
    x"0209000000000000015500000000000000fb33723f1c",
    x"030b0000000000000155fffffffffffff50003e7a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc93e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cfb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23b61c",
    x"070a0000000000000155fffffffffffff8ef35f92d1c",
    x"08020000000000000155fffffffffffff6f669e3021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a61c",
    x"0209000000000000015500000000000000fb3372391c",
    x"030b0000000000000155fffffffffffff50003e7a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc93c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cf71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23b01c",
    x"070a0000000000000155fffffffffffff8ef35f92a1c",
    x"08020000000000000155fffffffffffff6f669e3001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d29c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a71c",
    x"0209000000000000015500000000000000fb3372341c",
    x"030b0000000000000155fffffffffffff50003e7aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cf31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23a91c",
    x"070a0000000000000155fffffffffffff8ef35f9261c",
    x"08020000000000000155fffffffffffff6f669e2fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a81c",
    x"0209000000000000015500000000000000fb33722e1c",
    x"030b0000000000000155fffffffffffff50003e7ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cf01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23a31c",
    x"070a0000000000000155fffffffffffff8ef35f9221c",
    x"08020000000000000155fffffffffffff6f669e2fb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9a91c",
    x"0209000000000000015500000000000000fb3372291c",
    x"030b0000000000000155fffffffffffff50003e7ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd239d1c",
    x"070a0000000000000155fffffffffffff8ef35f91f1c",
    x"08020000000000000155fffffffffffff6f669e2f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9aa1c",
    x"0209000000000000015500000000000000fb3372231c",
    x"030b0000000000000155fffffffffffff50003e7ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ce81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23971c",
    x"070a0000000000000155fffffffffffff8ef35f91b1c",
    x"08020000000000000155fffffffffffff6f669e2f61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d28c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9ab1c",
    x"0209000000000000015500000000000000fb33721d1c",
    x"030b0000000000000155fffffffffffff50003e7ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc92f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ce51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23911c",
    x"070a0000000000000155fffffffffffff8ef35f9171c",
    x"08020000000000000155fffffffffffff6f669e2f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9ac1c",
    x"0209000000000000015500000000000000fb3372181c",
    x"030b0000000000000155fffffffffffff50003e7af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc92d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ce11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd238b1c",
    x"070a0000000000000155fffffffffffff8ef35f9141c",
    x"08020000000000000155fffffffffffff6f669e2f11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9ae1c",
    x"0209000000000000015500000000000000fb3372121c",
    x"030b0000000000000155fffffffffffff50003e7b01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc92b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cdd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23841c",
    x"070a0000000000000155fffffffffffff8ef35f9101c",
    x"08020000000000000155fffffffffffff6f669e2ef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d27f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9af1c",
    x"0209000000000000015500000000000000fb33720d1c",
    x"030b0000000000000155fffffffffffff50003e7b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cda1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd237e1c",
    x"070a0000000000000155fffffffffffff8ef35f90d1c",
    x"08020000000000000155fffffffffffff6f669e2ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d27b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9b01c",
    x"0209000000000000015500000000000000fb3372071c",
    x"030b0000000000000155fffffffffffff50003e7b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cd61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23781c",
    x"070a0000000000000155fffffffffffff8ef35f9091c",
    x"08020000000000000155fffffffffffff6f669e2ea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9b11c",
    x"0209000000000000015500000000000000fb3372011c",
    x"030b0000000000000155fffffffffffff50003e7b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cd31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23721c",
    x"070a0000000000000155fffffffffffff8ef35f9051c",
    x"08020000000000000155fffffffffffff6f669e2e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9b21c",
    x"0209000000000000015500000000000000fb3371fc1c",
    x"030b0000000000000155fffffffffffff50003e7b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ccf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd236c1c",
    x"070a0000000000000155fffffffffffff8ef35f9021c",
    x"08020000000000000155fffffffffffff6f669e2e51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d26e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9b31c",
    x"0209000000000000015500000000000000fb3371f61c",
    x"030b0000000000000155fffffffffffff50003e7b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc91e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ccb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23661c",
    x"070a0000000000000155fffffffffffff8ef35f8fe1c",
    x"08020000000000000155fffffffffffff6f669e2e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d26a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9b41c",
    x"0209000000000000031f00000000000000fb3371f11c",
    x"030b000000000000031ffffffffffffff50003e7b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc91c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3cc81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd23601c",
    x"070a000000000000031ffffffffffffff8ef35f8fa1c",
    x"0802000000000000031ffffffffffffff6f669e2e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d2661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9b51c",
    x"020900000000000000ae00000000000000fb3371eb1c",
    x"030b00000000000000aefffffffffffff50003e7b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc9191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3cc41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd23591c",
    x"070a00000000000000aefffffffffffff8ef35f8f71c",
    x"080200000000000000aefffffffffffff6f669e2de1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d2621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9b61c",
    x"020900000000000001a400000000000000fb3371e51c",
    x"030b00000000000001a4fffffffffffff50003e7b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc9171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3cc01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd23531c",
    x"070a00000000000001a4fffffffffffff8ef35f8f31c",
    x"080200000000000001a4fffffffffffff6f669e2dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266d25e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbe9b81c",
    x"0209000000000000015600000000000000fb3371e01c",
    x"030b0000000000000156fffffffffffff50003e7b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc9151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3cbd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd234d1c",
    x"070a0000000000000156fffffffffffff8ef35f8ef1c",
    x"08020000000000000156fffffffffffff6f669e2d91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d25a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9b91c",
    x"0209000000000000015500000000000000fb3371da1c",
    x"030b0000000000000155fffffffffffff50003e7ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cb91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23471c",
    x"070a0000000000000155fffffffffffff8ef35f8ec1c",
    x"08020000000000000155fffffffffffff6f669e2d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d2551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe9ba1c",
    x"0209000000000000016a00000000000000fb3371d51c",
    x"030b000000000000016afffffffffffff50003e7bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc9101c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3cb51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd23411c",
    x"070a000000000000016afffffffffffff8ef35f8e81c",
    x"0802000000000000016afffffffffffff6f669e2d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9bb1c",
    x"0209000000000000015500000000000000fb3371cf1c",
    x"030b0000000000000155fffffffffffff50003e7bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc90d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cb21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd233b1c",
    x"070a0000000000000155fffffffffffff8ef35f8e41c",
    x"08020000000000000155fffffffffffff6f669e2d21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d24d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9bc1c",
    x"0209000000000000015500000000000000fb3371c91c",
    x"030b0000000000000155fffffffffffff50003e7bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc90b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3cae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23341c",
    x"070a0000000000000155fffffffffffff8ef35f8e11c",
    x"08020000000000000155fffffffffffff6f669e2d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2491c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9bd1c",
    x"0209000000000000015500000000000000fb3371c41c",
    x"030b0000000000000155fffffffffffff50003e7be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3caa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd232e1c",
    x"070a0000000000000155fffffffffffff8ef35f8dd1c",
    x"08020000000000000155fffffffffffff6f669e2cd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2451c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9be1c",
    x"0209000000000000015500000000000000fb3371be1c",
    x"030b0000000000000155fffffffffffff50003e7be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9061c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ca71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23281c",
    x"070a0000000000000155fffffffffffff8ef35f8d91c",
    x"08020000000000000155fffffffffffff6f669e2cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9bf1c",
    x"0209000000000000015500000000000000fb3371b91c",
    x"030b0000000000000155fffffffffffff50003e7bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3ca31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23221c",
    x"070a0000000000000155fffffffffffff8ef35f8d61c",
    x"08020000000000000155fffffffffffff6f669e2c91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d23c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c11c",
    x"0209000000000000015500000000000000fb3371b31c",
    x"030b0000000000000155fffffffffffff50003e7c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc9011c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c9f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd231c1c",
    x"070a0000000000000155fffffffffffff8ef35f8d21c",
    x"08020000000000000155fffffffffffff6f669e2c61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c21c",
    x"0209000000000000015500000000000000fb3371ad1c",
    x"030b0000000000000155fffffffffffff50003e7c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8fe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c9c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23161c",
    x"070a0000000000000155fffffffffffff8ef35f8ce1c",
    x"08020000000000000155fffffffffffff6f669e2c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c31c",
    x"0209000000000000015500000000000000fb3371a81c",
    x"030b0000000000000155fffffffffffff50003e7c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8fc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd230f1c",
    x"070a0000000000000155fffffffffffff8ef35f8cb1c",
    x"08020000000000000155fffffffffffff6f669e2c11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c41c",
    x"0209000000000000015500000000000000fb3371a21c",
    x"030b0000000000000155fffffffffffff50003e7c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8fa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23091c",
    x"070a0000000000000155fffffffffffff8ef35f8c71c",
    x"08020000000000000155fffffffffffff6f669e2bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d22c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c51c",
    x"0209000000000000015500000000000000fb33719d1c",
    x"030b0000000000000155fffffffffffff50003e7c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8f71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd23031c",
    x"070a0000000000000155fffffffffffff8ef35f8c31c",
    x"08020000000000000155fffffffffffff6f669e2bd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c61c",
    x"0209000000000000015500000000000000fb3371971c",
    x"030b0000000000000155fffffffffffff50003e7c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8f51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c8d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd22fd1c",
    x"070a0000000000000155fffffffffffff8ef35f8c01c",
    x"08020000000000000155fffffffffffff6f669e2ba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d2231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c71c",
    x"0209000000000000015500000000000000fb3371911c",
    x"030b0000000000000155fffffffffffff50003e7c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8f21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd22f71c",
    x"070a0000000000000155fffffffffffff8ef35f8bc1c",
    x"08020000000000000155fffffffffffff6f669e2b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266d21f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a50000000000000b0bfbe9c81c",
    x"020900000000000001a500000000000000fb33718c1c",
    x"030b00000000000001a5fffffffffffff50003e7c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc8f01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f3c861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd22f11c",
    x"070a00000000000001a5fffffffffffff8ef35f8b91c",
    x"080200000000000001a5fffffffffffff6f669e2b51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d21b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9c91c",
    x"0209000000000000015500000000000000fb3371861c",
    x"030b0000000000000155fffffffffffff50003e7c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8ed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3c821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd22ea1c",
    x"070a0000000000000155fffffffffffff8ef35f8b51c",
    x"08020000000000000155fffffffffffff6f669e2b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d2171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9cb1c",
    x"0209000000000000031f00000000000000fb3371801c",
    x"030b000000000000031ffffffffffffff50003e7c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc8eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3c7e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd22e41c",
    x"070a000000000000031ffffffffffffff8ef35f8b11c",
    x"0802000000000000031ffffffffffffff6f669e2b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d2121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9cc1c",
    x"020900000000000000ae00000000000000fb33717b1c",
    x"030b00000000000000aefffffffffffff50003e7ca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc8e81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3c7b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd22de1c",
    x"070a00000000000000aefffffffffffff8ef35f8ae1c",
    x"080200000000000000aefffffffffffff6f669e2ae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d20e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9cd1c",
    x"020900000000000001a400000000000000fb3371751c",
    x"030b00000000000001a4fffffffffffff50003e7cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc8e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3c771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd22d81c",
    x"070a00000000000001a4fffffffffffff8ef35f8aa1c",
    x"080200000000000001a4fffffffffffff6f669e2ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266d20a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbe9ce1c",
    x"0209000000000000025600000000000000fb3371701c",
    x"030b0000000000000256fffffffffffff50003e7cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dc8e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f3c731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd22d21c",
    x"070a0000000000000256fffffffffffff8ef35f8a61c",
    x"08020000000000000256fffffffffffff6f669e2a91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d2061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9cf1c",
    x"020900000000000002aa00000000000000fb33716a1c",
    x"030b00000000000002aafffffffffffff50003e7cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c701c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22cc1c",
    x"070a00000000000002aafffffffffffff8ef35f8a31c",
    x"080200000000000002aafffffffffffff6f669e2a71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d2021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d01c",
    x"020900000000000002aa00000000000000fb3371641c",
    x"030b00000000000002aafffffffffffff50003e7ce1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c6c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22c51c",
    x"070a00000000000002aafffffffffffff8ef35f89f1c",
    x"080200000000000002aafffffffffffff6f669e2a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1fe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d11c",
    x"020900000000000002aa00000000000000fb33715f1c",
    x"030b00000000000002aafffffffffffff50003e7cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8dc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22bf1c",
    x"070a00000000000002aafffffffffffff8ef35f89b1c",
    x"080200000000000002aafffffffffffff6f669e2a21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d21c",
    x"020900000000000002aa00000000000000fb3371591c",
    x"030b00000000000002aafffffffffffff50003e7d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22b91c",
    x"070a00000000000002aafffffffffffff8ef35f8981c",
    x"080200000000000002aafffffffffffff6f669e2a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d41c",
    x"020900000000000002aa00000000000000fb3371541c",
    x"030b00000000000002aafffffffffffff50003e7d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8d71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22b31c",
    x"070a00000000000002aafffffffffffff8ef35f8941c",
    x"080200000000000002aafffffffffffff6f669e29d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1f11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d51c",
    x"020900000000000002aa00000000000000fb33714e1c",
    x"030b00000000000002aafffffffffffff50003e7d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8d51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c5d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22ad1c",
    x"070a00000000000002aafffffffffffff8ef35f8901c",
    x"080200000000000002aafffffffffffff6f669e29b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1ed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d61c",
    x"020900000000000002aa00000000000000fb3371481c",
    x"030b00000000000002aafffffffffffff50003e7d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8d21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c5a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22a71c",
    x"070a00000000000002aafffffffffffff8ef35f88d1c",
    x"080200000000000002aafffffffffffff6f669e2991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1e91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d71c",
    x"020900000000000002aa00000000000000fb3371431c",
    x"030b00000000000002aafffffffffffff50003e7d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8d01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22a01c",
    x"070a00000000000002aafffffffffffff8ef35f8891c",
    x"080200000000000002aafffffffffffff6f669e2961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d81c",
    x"020900000000000002aa00000000000000fb33713d1c",
    x"030b00000000000002aafffffffffffff50003e7d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8ce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd229a1c",
    x"070a00000000000002aafffffffffffff8ef35f8851c",
    x"080200000000000002aafffffffffffff6f669e2941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9d91c",
    x"020900000000000002aa00000000000000fb3371381c",
    x"030b00000000000002aafffffffffffff50003e7d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8cb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c4f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22941c",
    x"070a00000000000002aafffffffffffff8ef35f8821c",
    x"080200000000000002aafffffffffffff6f669e2911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1dc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9da1c",
    x"020900000000000002aa00000000000000fb3371321c",
    x"030b00000000000002aafffffffffffff50003e7d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8c91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c4b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd228e1c",
    x"070a00000000000002aafffffffffffff8ef35f87e1c",
    x"080200000000000002aafffffffffffff6f669e28f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9db1c",
    x"020900000000000002aa00000000000000fb33712c1c",
    x"030b00000000000002aafffffffffffff50003e7d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8c61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22881c",
    x"070a00000000000002aafffffffffffff8ef35f87a1c",
    x"080200000000000002aafffffffffffff6f669e28d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1d41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9dc1c",
    x"020900000000000002aa00000000000000fb3371271c",
    x"030b00000000000002aafffffffffffff50003e7d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8c41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22821c",
    x"070a00000000000002aafffffffffffff8ef35f8771c",
    x"080200000000000002aafffffffffffff6f669e28a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1d01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9de1c",
    x"020900000000000002aa00000000000000fb3371211c",
    x"030b00000000000002aafffffffffffff50003e7d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8c11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd227c1c",
    x"070a00000000000002aafffffffffffff8ef35f8731c",
    x"080200000000000002aafffffffffffff6f669e2881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266d1cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbe9df1c",
    x"0209000000000000029a00000000000000fb33711c1c",
    x"030b000000000000029afffffffffffff50003e7da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc8bf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f3c3d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd22751c",
    x"070a000000000000029afffffffffffff8ef35f86f1c",
    x"0802000000000000029afffffffffffff6f669e2851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9e01c",
    x"020900000000000002aa00000000000000fb3371161c",
    x"030b00000000000002aafffffffffffff50003e7db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8bc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd226f1c",
    x"070a00000000000002aafffffffffffff8ef35f86c1c",
    x"080200000000000002aafffffffffffff6f669e2831c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d1c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9e11c",
    x"0209000000000000031f00000000000000fb3371101c",
    x"030b000000000000031ffffffffffffff50003e7dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc8ba1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3c351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd22691c",
    x"070a000000000000031ffffffffffffff8ef35f8681c",
    x"0802000000000000031ffffffffffffff6f669e2811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d1bf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9e21c",
    x"020900000000000000ae00000000000000fb33710b1c",
    x"030b00000000000000aefffffffffffff50003e7dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc8b71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3c321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd22631c",
    x"070a00000000000000aefffffffffffff8ef35f8651c",
    x"080200000000000000aefffffffffffff6f669e27e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d1bb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9e31c",
    x"020900000000000001a400000000000000fb3371051c",
    x"030b00000000000001a4fffffffffffff50003e7de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc8b51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3c2e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd225d1c",
    x"070a00000000000001a4fffffffffffff8ef35f8611c",
    x"080200000000000001a4fffffffffffff6f669e27c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266d1b71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbe9e41c",
    x"0209000000000000029600000000000000fb3371001c",
    x"030b0000000000000296fffffffffffff50003e7df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dc8b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f3c2a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd22571c",
    x"070a0000000000000296fffffffffffff8ef35f85d1c",
    x"08020000000000000296fffffffffffff6f669e2791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266d1b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbe9e51c",
    x"0209000000000000016a00000000000000fb3370fa1c",
    x"030b000000000000016afffffffffffff50003e7e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc8b01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3c271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd22501c",
    x"070a000000000000016afffffffffffff8ef35f85a1c",
    x"0802000000000000016afffffffffffff6f669e2771c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000299ffffffffffffff0266d1ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002990000000000000b0bfbe9e61c",
    x"0209000000000000029900000000000000fb3370f41c",
    x"030b0000000000000299fffffffffffff50003e7e11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc8ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002990000000000000b072f3c231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002990000000000000004cd224a1c",
    x"070a0000000000000299fffffffffffff8ef35f8561c",
    x"08020000000000000299fffffffffffff6f669e2751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9e81c",
    x"020900000000000002aa00000000000000fb3370ef1c",
    x"030b00000000000002aafffffffffffff50003e7e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8ab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c1f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22441c",
    x"070a00000000000002aafffffffffffff8ef35f8521c",
    x"080200000000000002aafffffffffffff6f669e2721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1a61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9e91c",
    x"020900000000000002aa00000000000000fb3370e91c",
    x"030b00000000000002aafffffffffffff50003e7e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c1c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd223e1c",
    x"070a00000000000002aafffffffffffff8ef35f84f1c",
    x"080200000000000002aafffffffffffff6f669e2701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9ea1c",
    x"020900000000000002aa00000000000000fb3370e41c",
    x"030b00000000000002aafffffffffffff50003e7e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8a61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22381c",
    x"070a00000000000002aafffffffffffff8ef35f84b1c",
    x"080200000000000002aafffffffffffff6f669e26d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d19d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9eb1c",
    x"020900000000000002aa00000000000000fb3370de1c",
    x"030b00000000000002aafffffffffffff50003e7e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22321c",
    x"070a00000000000002aafffffffffffff8ef35f8471c",
    x"080200000000000002aafffffffffffff6f669e26b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9ec1c",
    x"020900000000000002aa00000000000000fb3370d81c",
    x"030b00000000000002aafffffffffffff50003e7e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8a11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd222b1c",
    x"070a00000000000002aafffffffffffff8ef35f8441c",
    x"080200000000000002aafffffffffffff6f669e2691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9ed1c",
    x"020900000000000002aa00000000000000fb3370d31c",
    x"030b00000000000002aafffffffffffff50003e7e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc89f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c0d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22251c",
    x"070a00000000000002aafffffffffffff8ef35f8401c",
    x"080200000000000002aafffffffffffff6f669e2661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9ee1c",
    x"020900000000000002aa00000000000000fb3370cd1c",
    x"030b00000000000002aafffffffffffff50003e7e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc89d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd221f1c",
    x"070a00000000000002aafffffffffffff8ef35f83c1c",
    x"080200000000000002aafffffffffffff6f669e2641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d18d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9ef1c",
    x"020900000000000002aa00000000000000fb3370c71c",
    x"030b00000000000002aafffffffffffff50003e7e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc89a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22191c",
    x"070a00000000000002aafffffffffffff8ef35f8391c",
    x"080200000000000002aafffffffffffff6f669e2611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1891c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9f11c",
    x"020900000000000002aa00000000000000fb3370c21c",
    x"030b00000000000002aafffffffffffff50003e7e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3c021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22131c",
    x"070a00000000000002aafffffffffffff8ef35f8351c",
    x"080200000000000002aafffffffffffff6f669e25f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9f21c",
    x"020900000000000002aa00000000000000fb3370bc1c",
    x"030b00000000000002aafffffffffffff50003e7ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3bfe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd220d1c",
    x"070a00000000000002aafffffffffffff8ef35f8311c",
    x"080200000000000002aafffffffffffff6f669e25d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9f31c",
    x"020900000000000002aa00000000000000fb3370b71c",
    x"030b00000000000002aafffffffffffff50003e7eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3bfb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22061c",
    x"070a00000000000002aafffffffffffff8ef35f82e1c",
    x"080200000000000002aafffffffffffff6f669e25a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d17c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9f41c",
    x"020900000000000002aa00000000000000fb3370b11c",
    x"030b00000000000002aafffffffffffff50003e7ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3bf71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd22001c",
    x"070a00000000000002aafffffffffffff8ef35f82a1c",
    x"080200000000000002aafffffffffffff6f669e2581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbe9f51c",
    x"020900000000000002aa00000000000000fb3370ab1c",
    x"030b00000000000002aafffffffffffff50003e7ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc88e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3bf31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21fa1c",
    x"070a00000000000002aafffffffffffff8ef35f8261c",
    x"080200000000000002aafffffffffffff6f669e2551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1741c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9f61c",
    x"0209000000000000015500000000000000fb3370a61c",
    x"030b0000000000000155fffffffffffff50003e7ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc88b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bf01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21f41c",
    x"070a0000000000000155fffffffffffff8ef35f8231c",
    x"08020000000000000155fffffffffffff6f669e2531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d16f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbe9f71c",
    x"0209000000000000031f00000000000000fb3370a01c",
    x"030b000000000000031ffffffffffffff50003e7ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc8891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3bec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd21ee1c",
    x"070a000000000000031ffffffffffffff8ef35f81f1c",
    x"0802000000000000031ffffffffffffff6f669e2511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d16b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbe9f81c",
    x"020900000000000000ae00000000000000fb33709b1c",
    x"030b00000000000000aefffffffffffff50003e7f01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc8861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3be91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd21e81c",
    x"070a00000000000000aefffffffffffff8ef35f81b1c",
    x"080200000000000000aefffffffffffff6f669e24e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d1671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbe9fa1c",
    x"020900000000000001a400000000000000fb3370951c",
    x"030b00000000000001a4fffffffffffff50003e7f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc8841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3be51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd21e11c",
    x"070a00000000000001a4fffffffffffff8ef35f8181c",
    x"080200000000000001a4fffffffffffff6f669e24c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266d1631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbe9fb1c",
    x"0209000000000000019600000000000000fb33708f1c",
    x"030b0000000000000196fffffffffffff50003e7f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc8821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f3be11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001960000000000000004cd21db1c",
    x"070a0000000000000196fffffffffffff8ef35f8141c",
    x"08020000000000000196fffffffffffff6f669e2491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d15f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9fc1c",
    x"0209000000000000015500000000000000fb33708a1c",
    x"030b0000000000000155fffffffffffff50003e7f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc87f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bde1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21d51c",
    x"070a0000000000000155fffffffffffff8ef35f8101c",
    x"08020000000000000155fffffffffffff6f669e2471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d15b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9fd1c",
    x"0209000000000000015500000000000000fb3370841c",
    x"030b0000000000000155fffffffffffff50003e7f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc87d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bda1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21cf1c",
    x"070a0000000000000155fffffffffffff8ef35f80d1c",
    x"08020000000000000155fffffffffffff6f669e2451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9fe1c",
    x"0209000000000000015500000000000000fb33707f1c",
    x"030b0000000000000155fffffffffffff50003e7f51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc87a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bd61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21c91c",
    x"070a0000000000000155fffffffffffff8ef35f8091c",
    x"08020000000000000155fffffffffffff6f669e2421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbe9ff1c",
    x"0209000000000000015500000000000000fb3370791c",
    x"030b0000000000000155fffffffffffff50003e7f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bd31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21c31c",
    x"070a0000000000000155fffffffffffff8ef35f8051c",
    x"08020000000000000155fffffffffffff6f669e2401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d14e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea001c",
    x"0209000000000000015500000000000000fb3370731c",
    x"030b0000000000000155fffffffffffff50003e7f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bcf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21bc1c",
    x"070a0000000000000155fffffffffffff8ef35f8021c",
    x"08020000000000000155fffffffffffff6f669e23d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d14a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea011c",
    x"0209000000000000015500000000000000fb33706e1c",
    x"030b0000000000000155fffffffffffff50003e7f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bcb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21b61c",
    x"070a0000000000000155fffffffffffff8ef35f7fe1c",
    x"08020000000000000155fffffffffffff6f669e23b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea021c",
    x"0209000000000000015500000000000000fb3370681c",
    x"030b0000000000000155fffffffffffff50003e7f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bc81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21b01c",
    x"070a0000000000000155fffffffffffff8ef35f7fa1c",
    x"08020000000000000155fffffffffffff6f669e2391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea041c",
    x"0209000000000000015500000000000000fb3370631c",
    x"030b0000000000000155fffffffffffff50003e7fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc86e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bc41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21aa1c",
    x"070a0000000000000155fffffffffffff8ef35f7f71c",
    x"08020000000000000155fffffffffffff6f669e2361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d13d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea051c",
    x"0209000000000000015500000000000000fb33705d1c",
    x"030b0000000000000155fffffffffffff50003e7fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc86b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bc01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21a41c",
    x"070a0000000000000155fffffffffffff8ef35f7f31c",
    x"08020000000000000155fffffffffffff6f669e2341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea061c",
    x"0209000000000000015500000000000000fb3370571c",
    x"030b0000000000000155fffffffffffff50003e7fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bbd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd219e1c",
    x"070a0000000000000155fffffffffffff8ef35f7f01c",
    x"08020000000000000155fffffffffffff6f669e2311c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea071c",
    x"0209000000000000015500000000000000fb3370521c",
    x"030b0000000000000155fffffffffffff50003e7fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bb91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21971c",
    x"070a0000000000000155fffffffffffff8ef35f7ec1c",
    x"08020000000000000155fffffffffffff6f669e22f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea081c",
    x"0209000000000000015500000000000000fb33704c1c",
    x"030b0000000000000155fffffffffffff50003e7fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bb51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21911c",
    x"070a0000000000000155fffffffffffff8ef35f7e81c",
    x"08020000000000000155fffffffffffff6f669e22d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d12d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea091c",
    x"0209000000000000015500000000000000fb3370471c",
    x"030b0000000000000155fffffffffffff50003e7fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8621c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bb21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd218b1c",
    x"070a0000000000000155fffffffffffff8ef35f7e51c",
    x"08020000000000000155fffffffffffff6f669e22a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d1281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea0a1c",
    x"0209000000000000015500000000000000fb3370411c",
    x"030b0000000000000155fffffffffffff50003e7ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc85f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3bae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd21851c",
    x"070a0000000000000155fffffffffffff8ef35f7e11c",
    x"08020000000000000155fffffffffffff6f669e2281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266d1241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbea0b1c",
    x"020900000000000002a500000000000000fb33703b1c",
    x"030b00000000000002a5fffffffffffff50003e8001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc85d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f3baa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd217f1c",
    x"070a00000000000002a5fffffffffffff8ef35f7dd1c",
    x"080200000000000002a5fffffffffffff6f669e2251c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea0d1c",
    x"020900000000000002aa00000000000000fb3370361c",
    x"030b00000000000002aafffffffffffff50003e8011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc85a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ba71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21791c",
    x"070a00000000000002aafffffffffffff8ef35f7da1c",
    x"080200000000000002aafffffffffffff6f669e2231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d11c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea0e1c",
    x"0209000000000000031f00000000000000fb3370301c",
    x"030b000000000000031ffffffffffffff50003e8021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc8581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3ba31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd21731c",
    x"070a000000000000031ffffffffffffff8ef35f7d61c",
    x"0802000000000000031ffffffffffffff6f669e2211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d1181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea0f1c",
    x"020900000000000000ae00000000000000fb33702a1c",
    x"030b00000000000000aefffffffffffff50003e8031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc8551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3b9f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd216c1c",
    x"070a00000000000000aefffffffffffff8ef35f7d21c",
    x"080200000000000000aefffffffffffff6f669e21e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d1141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea101c",
    x"020900000000000001a400000000000000fb3370251c",
    x"030b00000000000001a4fffffffffffff50003e8041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc8531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3b9c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd21661c",
    x"070a00000000000001a4fffffffffffff8ef35f7cf1c",
    x"080200000000000001a4fffffffffffff6f669e21c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d10f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbea111c",
    x"020900000000000002a600000000000000fb33701f1c",
    x"030b00000000000002a6fffffffffffff50003e8051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc8501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3b981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd21601c",
    x"070a00000000000002a6fffffffffffff8ef35f7cb1c",
    x"080200000000000002a6fffffffffffff6f669e2191c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d10b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea121c",
    x"020900000000000002aa00000000000000fb33701a1c",
    x"030b00000000000002aafffffffffffff50003e8061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc84e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd215a1c",
    x"070a00000000000002aafffffffffffff8ef35f7c71c",
    x"080200000000000002aafffffffffffff6f669e2171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266d1071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbea131c",
    x"020900000000000002a600000000000000fb3370141c",
    x"030b00000000000002a6fffffffffffff50003e8071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc84c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3b911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd21541c",
    x"070a00000000000002a6fffffffffffff8ef35f7c41c",
    x"080200000000000002a6fffffffffffff6f669e2151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d1031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea141c",
    x"020900000000000002aa00000000000000fb33700e1c",
    x"030b00000000000002aafffffffffffff50003e8081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b8d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd214e1c",
    x"070a00000000000002aafffffffffffff8ef35f7c01c",
    x"080200000000000002aafffffffffffff6f669e2121c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea151c",
    x"020900000000000002aa00000000000000fb3370091c",
    x"030b00000000000002aafffffffffffff50003e8091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b8a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21471c",
    x"070a00000000000002aafffffffffffff8ef35f7bc1c",
    x"080200000000000002aafffffffffffff6f669e2101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0fa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea171c",
    x"020900000000000002aa00000000000000fb3370031c",
    x"030b00000000000002aafffffffffffff50003e80a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21411c",
    x"070a00000000000002aafffffffffffff8ef35f7b91c",
    x"080200000000000002aafffffffffffff6f669e20d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0f61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea181c",
    x"020900000000000002aa00000000000000fb336ffe1c",
    x"030b00000000000002aafffffffffffff50003e80b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd213b1c",
    x"070a00000000000002aafffffffffffff8ef35f7b51c",
    x"080200000000000002aafffffffffffff6f669e20b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0f21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea191c",
    x"020900000000000002aa00000000000000fb336ff81c",
    x"030b00000000000002aafffffffffffff50003e80c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc83f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b7f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21351c",
    x"070a00000000000002aafffffffffffff8ef35f7b11c",
    x"080200000000000002aafffffffffffff6f669e2091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea1a1c",
    x"020900000000000002aa00000000000000fb336ff21c",
    x"030b00000000000002aafffffffffffff50003e80d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc83d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b7b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd212f1c",
    x"070a00000000000002aafffffffffffff8ef35f7ae1c",
    x"080200000000000002aafffffffffffff6f669e2061c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0ea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea1b1c",
    x"020900000000000002aa00000000000000fb336fed1c",
    x"030b00000000000002aafffffffffffff50003e80e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc83a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21291c",
    x"070a00000000000002aafffffffffffff8ef35f7aa1c",
    x"080200000000000002aafffffffffffff6f669e2041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0e61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea1c1c",
    x"020900000000000002aa00000000000000fb336fe71c",
    x"030b00000000000002aafffffffffffff50003e80e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21221c",
    x"070a00000000000002aafffffffffffff8ef35f7a61c",
    x"080200000000000002aafffffffffffff6f669e2011c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0e11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea1d1c",
    x"020900000000000002aa00000000000000fb336fe21c",
    x"030b00000000000002aafffffffffffff50003e80f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8351c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b701c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd211c1c",
    x"070a00000000000002aafffffffffffff8ef35f7a31c",
    x"080200000000000002aafffffffffffff6f669e1ff1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0dd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea1e1c",
    x"020900000000000002aa00000000000000fb336fdc1c",
    x"030b00000000000002aafffffffffffff50003e8101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b6c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21161c",
    x"070a00000000000002aafffffffffffff8ef35f79f1c",
    x"080200000000000002aafffffffffffff6f669e1fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0d91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea201c",
    x"020900000000000002aa00000000000000fb336fd61c",
    x"030b00000000000002aafffffffffffff50003e8111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21101c",
    x"070a00000000000002aafffffffffffff8ef35f79b1c",
    x"080200000000000002aafffffffffffff6f669e1fa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0d51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea211c",
    x"020900000000000002aa00000000000000fb336fd11c",
    x"030b00000000000002aafffffffffffff50003e8121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc82e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd210a1c",
    x"070a00000000000002aafffffffffffff8ef35f7981c",
    x"080200000000000002aafffffffffffff6f669e1f81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0d11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea221c",
    x"020900000000000002aa00000000000000fb336fcb1c",
    x"030b00000000000002aafffffffffffff50003e8131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc82c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd21041c",
    x"070a00000000000002aafffffffffffff8ef35f7941c",
    x"080200000000000002aafffffffffffff6f669e1f51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0cd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea231c",
    x"020900000000000002aa00000000000000fb336fc61c",
    x"030b00000000000002aafffffffffffff50003e8141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc8291c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b5e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20fd1c",
    x"070a00000000000002aafffffffffffff8ef35f7901c",
    x"080200000000000002aafffffffffffff6f669e1f31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d0c81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea241c",
    x"0209000000000000031f00000000000000fb336fc01c",
    x"030b000000000000031ffffffffffffff50003e8151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc8271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3b5a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd20f71c",
    x"070a000000000000031ffffffffffffff8ef35f78d1c",
    x"0802000000000000031ffffffffffffff6f669e1f11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d0c41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea251c",
    x"020900000000000000ae00000000000000fb336fba1c",
    x"030b00000000000000aefffffffffffff50003e8161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc8241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3b561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd20f11c",
    x"070a00000000000000aefffffffffffff8ef35f7891c",
    x"080200000000000000aefffffffffffff6f669e1ee1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d0c01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea261c",
    x"020900000000000001a400000000000000fb336fb51c",
    x"030b00000000000001a4fffffffffffff50003e8171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc8221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3b531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd20eb1c",
    x"070a00000000000001a4fffffffffffff8ef35f7851c",
    x"080200000000000001a4fffffffffffff6f669e1ec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266d0bc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbea271c",
    x"020900000000000001a600000000000000fb336faf1c",
    x"030b00000000000001a6fffffffffffff50003e8181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc81f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f3b4f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd20e51c",
    x"070a00000000000001a6fffffffffffff8ef35f7821c",
    x"080200000000000001a6fffffffffffff6f669e1e91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0b81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea281c",
    x"0209000000000000015500000000000000fb336faa1c",
    x"030b0000000000000155fffffffffffff50003e8191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc81d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b4b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20df1c",
    x"070a0000000000000155fffffffffffff8ef35f77e1c",
    x"08020000000000000155fffffffffffff6f669e1e71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0b31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea2a1c",
    x"0209000000000000015500000000000000fb336fa41c",
    x"030b0000000000000155fffffffffffff50003e81a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc81a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20d81c",
    x"070a0000000000000155fffffffffffff8ef35f77a1c",
    x"08020000000000000155fffffffffffff6f669e1e51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0af1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea2b1c",
    x"0209000000000000015500000000000000fb336f9e1c",
    x"030b0000000000000155fffffffffffff50003e81b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20d21c",
    x"070a0000000000000155fffffffffffff8ef35f7771c",
    x"08020000000000000155fffffffffffff6f669e1e21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0ab1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea2c1c",
    x"0209000000000000015500000000000000fb336f991c",
    x"030b0000000000000155fffffffffffff50003e81c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20cc1c",
    x"070a0000000000000155fffffffffffff8ef35f7731c",
    x"08020000000000000155fffffffffffff6f669e1e01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0a71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea2d1c",
    x"0209000000000000015500000000000000fb336f931c",
    x"030b0000000000000155fffffffffffff50003e81d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b3d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20c61c",
    x"070a0000000000000155fffffffffffff8ef35f76f1c",
    x"08020000000000000155fffffffffffff6f669e1dd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0a31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea2e1c",
    x"0209000000000000015500000000000000fb336f8d1c",
    x"030b0000000000000155fffffffffffff50003e81e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20c01c",
    x"070a0000000000000155fffffffffffff8ef35f76c1c",
    x"08020000000000000155fffffffffffff6f669e1db1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d09f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea2f1c",
    x"0209000000000000015500000000000000fb336f881c",
    x"030b0000000000000155fffffffffffff50003e81f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc80e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20ba1c",
    x"070a0000000000000155fffffffffffff8ef35f7681c",
    x"08020000000000000155fffffffffffff6f669e1d91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d09a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea301c",
    x"0209000000000000015500000000000000fb336f821c",
    x"030b0000000000000155fffffffffffff50003e8201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc80c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20b31c",
    x"070a0000000000000155fffffffffffff8ef35f7641c",
    x"08020000000000000155fffffffffffff6f669e1d61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0961c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea311c",
    x"0209000000000000015500000000000000fb336f7d1c",
    x"030b0000000000000155fffffffffffff50003e8201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b2e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20ad1c",
    x"070a0000000000000155fffffffffffff8ef35f7611c",
    x"08020000000000000155fffffffffffff6f669e1d41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0921c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea331c",
    x"0209000000000000015500000000000000fb336f771c",
    x"030b0000000000000155fffffffffffff50003e8211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b2b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20a71c",
    x"070a0000000000000155fffffffffffff8ef35f75d1c",
    x"08020000000000000155fffffffffffff6f669e1d11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d08e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea341c",
    x"0209000000000000015500000000000000fb336f711c",
    x"030b0000000000000155fffffffffffff50003e8221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20a11c",
    x"070a0000000000000155fffffffffffff8ef35f7591c",
    x"08020000000000000155fffffffffffff6f669e1cf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d08a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea351c",
    x"0209000000000000015500000000000000fb336f6c1c",
    x"030b0000000000000155fffffffffffff50003e8231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc8021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd209b1c",
    x"070a0000000000000155fffffffffffff8ef35f7561c",
    x"08020000000000000155fffffffffffff6f669e1cd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0861c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea361c",
    x"0209000000000000015500000000000000fb336f661c",
    x"030b0000000000000155fffffffffffff50003e8241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc7ff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20951c",
    x"070a0000000000000155fffffffffffff8ef35f7521c",
    x"08020000000000000155fffffffffffff6f669e1ca1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0811c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea371c",
    x"0209000000000000015500000000000000fb336f611c",
    x"030b0000000000000155fffffffffffff50003e8251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc7fd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b1c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd208e1c",
    x"070a0000000000000155fffffffffffff8ef35f74e1c",
    x"08020000000000000155fffffffffffff6f669e1c81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266d07d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbea381c",
    x"0209000000000000029500000000000000fb336f5b1c",
    x"030b0000000000000295fffffffffffff50003e8261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc7fb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3b181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd20881c",
    x"070a0000000000000295fffffffffffff8ef35f74b1c",
    x"08020000000000000295fffffffffffff6f669e1c51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0791c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea391c",
    x"020900000000000002aa00000000000000fb336f551c",
    x"030b00000000000002aafffffffffffff50003e8271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3b151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20821c",
    x"070a00000000000002aafffffffffffff8ef35f7471c",
    x"080200000000000002aafffffffffffff6f669e1c31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d0751c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea3a1c",
    x"0209000000000000031f00000000000000fb336f501c",
    x"030b000000000000031ffffffffffffff50003e8281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc7f61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3b111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd207c1c",
    x"070a000000000000031ffffffffffffff8ef35f7431c",
    x"0802000000000000031ffffffffffffff6f669e1c11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d0711c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea3c1c",
    x"020900000000000000ae00000000000000fb336f4a1c",
    x"030b00000000000000aefffffffffffff50003e8291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc7f31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3b0d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd20761c",
    x"070a00000000000000aefffffffffffff8ef35f7401c",
    x"080200000000000000aefffffffffffff6f669e1be1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d06c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea3d1c",
    x"020900000000000001a400000000000000fb336f451c",
    x"030b00000000000001a4fffffffffffff50003e82a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc7f11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3b0a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd20701c",
    x"070a00000000000001a4fffffffffffff8ef35f73c1c",
    x"080200000000000001a4fffffffffffff6f669e1bc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266d0681c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbea3e1c",
    x"0209000000000000016600000000000000fb336f3f1c",
    x"030b0000000000000166fffffffffffff50003e82b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc7ee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f3b061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd20691c",
    x"070a0000000000000166fffffffffffff8ef35f7381c",
    x"08020000000000000166fffffffffffff6f669e1b91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266d0641c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea3f1c",
    x"0209000000000000015500000000000000fb336f391c",
    x"030b0000000000000155fffffffffffff50003e82c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc7ec1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3b021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd20631c",
    x"070a0000000000000155fffffffffffff8ef35f7351c",
    x"08020000000000000155fffffffffffff6f669e1b71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266d0601c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbea401c",
    x"020900000000000002a900000000000000fb336f341c",
    x"030b00000000000002a9fffffffffffff50003e82d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a9fffffffffffff4099dc7e91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f3aff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd205d1c",
    x"070a00000000000002a9fffffffffffff8ef35f7311c",
    x"080200000000000002a9fffffffffffff6f669e1b51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d05c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea411c",
    x"020900000000000002aa00000000000000fb336f2e1c",
    x"030b00000000000002aafffffffffffff50003e82e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7e71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3afb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20571c",
    x"070a00000000000002aafffffffffffff8ef35f72d1c",
    x"080200000000000002aafffffffffffff6f669e1b21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0581c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea421c",
    x"020900000000000002aa00000000000000fb336f291c",
    x"030b00000000000002aafffffffffffff50003e82f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3af81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20511c",
    x"070a00000000000002aafffffffffffff8ef35f72a1c",
    x"080200000000000002aafffffffffffff6f669e1b01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0531c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea431c",
    x"020900000000000002aa00000000000000fb336f231c",
    x"030b00000000000002aafffffffffffff50003e8301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7e21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3af41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd204b1c",
    x"070a00000000000002aafffffffffffff8ef35f7261c",
    x"080200000000000002aafffffffffffff6f669e1ad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d04f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea441c",
    x"020900000000000002aa00000000000000fb336f1d1c",
    x"030b00000000000002aafffffffffffff50003e8311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3af01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20441c",
    x"070a00000000000002aafffffffffffff8ef35f7221c",
    x"080200000000000002aafffffffffffff6f669e1ab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d04b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea461c",
    x"020900000000000002aa00000000000000fb336f181c",
    x"030b00000000000002aafffffffffffff50003e8311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7dd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd203e1c",
    x"070a00000000000002aafffffffffffff8ef35f71f1c",
    x"080200000000000002aafffffffffffff6f669e1a91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0471c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea471c",
    x"020900000000000002aa00000000000000fb336f121c",
    x"030b00000000000002aafffffffffffff50003e8321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7db1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ae91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20381c",
    x"070a00000000000002aafffffffffffff8ef35f71b1c",
    x"080200000000000002aafffffffffffff6f669e1a61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0431c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea481c",
    x"020900000000000002aa00000000000000fb336f0c1c",
    x"030b00000000000002aafffffffffffff50003e8331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7d81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ae51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20321c",
    x"070a00000000000002aafffffffffffff8ef35f7181c",
    x"080200000000000002aafffffffffffff6f669e1a41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d03f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea491c",
    x"020900000000000002aa00000000000000fb336f071c",
    x"030b00000000000002aafffffffffffff50003e8341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7d61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ae21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd202c1c",
    x"070a00000000000002aafffffffffffff8ef35f7141c",
    x"080200000000000002aafffffffffffff6f669e1a11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d03a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea4a1c",
    x"020900000000000002aa00000000000000fb336f011c",
    x"030b00000000000002aafffffffffffff50003e8351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7d31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ade1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20261c",
    x"070a00000000000002aafffffffffffff8ef35f7101c",
    x"080200000000000002aafffffffffffff6f669e19f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0361c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea4b1c",
    x"020900000000000002aa00000000000000fb336efc1c",
    x"030b00000000000002aafffffffffffff50003e8361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7d11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ada1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd201f1c",
    x"070a00000000000002aafffffffffffff8ef35f70d1c",
    x"080200000000000002aafffffffffffff6f669e19d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0321c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea4c1c",
    x"020900000000000002aa00000000000000fb336ef61c",
    x"030b00000000000002aafffffffffffff50003e8371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7ce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ad71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20191c",
    x"070a00000000000002aafffffffffffff8ef35f7091c",
    x"080200000000000002aafffffffffffff6f669e19a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d02e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea4d1c",
    x"020900000000000002aa00000000000000fb336ef01c",
    x"030b00000000000002aafffffffffffff50003e8381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ad31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20131c",
    x"070a00000000000002aafffffffffffff8ef35f7051c",
    x"080200000000000002aafffffffffffff6f669e1981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266d02a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbea4f1c",
    x"0209000000000000015a00000000000000fb336eeb1c",
    x"030b000000000000015afffffffffffff50003e8391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc7c91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3acf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd200d1c",
    x"070a000000000000015afffffffffffff8ef35f7021c",
    x"0802000000000000015afffffffffffff6f669e1951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0251c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea501c",
    x"020900000000000002aa00000000000000fb336ee51c",
    x"030b00000000000002aafffffffffffff50003e83a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3acc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd20071c",
    x"070a00000000000002aafffffffffffff8ef35f6fe1c",
    x"080200000000000002aafffffffffffff6f669e1931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266d0211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea511c",
    x"0209000000000000031f00000000000000fb336ee01c",
    x"030b000000000000031ffffffffffffff50003e83b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc7c41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3ac81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd20011c",
    x"070a000000000000031ffffffffffffff8ef35f6fa1c",
    x"0802000000000000031ffffffffffffff6f669e1911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266d01d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea521c",
    x"020900000000000000ae00000000000000fb336eda1c",
    x"030b00000000000000aefffffffffffff50003e83c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc7c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3ac41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1ffa1c",
    x"070a00000000000000aefffffffffffff8ef35f6f71c",
    x"080200000000000000aefffffffffffff6f669e18e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266d0191c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea531c",
    x"020900000000000001a400000000000000fb336ed41c",
    x"030b00000000000001a4fffffffffffff50003e83d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc7bf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3ac11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1ff41c",
    x"070a00000000000001a4fffffffffffff8ef35f6f31c",
    x"080200000000000001a4fffffffffffff6f669e18c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266d0151c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbea541c",
    x"0209000000000000026600000000000000fb336ecf1c",
    x"030b0000000000000266fffffffffffff50003e83e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc7bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f3abd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002660000000000000004cd1fee1c",
    x"070a0000000000000266fffffffffffff8ef35f6ef1c",
    x"08020000000000000266fffffffffffff6f669e1891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea551c",
    x"020900000000000002aa00000000000000fb336ec91c",
    x"030b00000000000002aafffffffffffff50003e83f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fe81c",
    x"070a00000000000002aafffffffffffff8ef35f6ec1c",
    x"080200000000000002aafffffffffffff6f669e1871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d00c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea561c",
    x"020900000000000002aa00000000000000fb336ec41c",
    x"030b00000000000002aafffffffffffff50003e8401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ab61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fe21c",
    x"070a00000000000002aafffffffffffff8ef35f6e81c",
    x"080200000000000002aafffffffffffff6f669e1851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0081c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea581c",
    x"020900000000000002aa00000000000000fb336ebe1c",
    x"030b00000000000002aafffffffffffff50003e8411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3ab21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fdc1c",
    x"070a00000000000002aafffffffffffff8ef35f6e41c",
    x"080200000000000002aafffffffffffff6f669e1821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0041c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea591c",
    x"020900000000000002aa00000000000000fb336eb81c",
    x"030b00000000000002aafffffffffffff50003e8421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aaf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fd51c",
    x"070a00000000000002aafffffffffffff8ef35f6e11c",
    x"080200000000000002aafffffffffffff6f669e1801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266d0001c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea5a1c",
    x"020900000000000002aa00000000000000fb336eb31c",
    x"030b00000000000002aafffffffffffff50003e8421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7b11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fcf1c",
    x"070a00000000000002aafffffffffffff8ef35f6dd1c",
    x"080200000000000002aafffffffffffff6f669e17d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cffc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea5b1c",
    x"020900000000000002aa00000000000000fb336ead1c",
    x"030b00000000000002aafffffffffffff50003e8431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aa71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fc91c",
    x"070a00000000000002aafffffffffffff8ef35f6d91c",
    x"080200000000000002aafffffffffffff6f669e17b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cff81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea5c1c",
    x"020900000000000002aa00000000000000fb336ea81c",
    x"030b00000000000002aafffffffffffff50003e8441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7ac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aa41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fc31c",
    x"070a00000000000002aafffffffffffff8ef35f6d61c",
    x"080200000000000002aafffffffffffff6f669e1791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cff31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea5d1c",
    x"020900000000000002aa00000000000000fb336ea21c",
    x"030b00000000000002aafffffffffffff50003e8451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3aa01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fbd1c",
    x"070a00000000000002aafffffffffffff8ef35f6d21c",
    x"080200000000000002aafffffffffffff6f669e1761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfef1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea5e1c",
    x"020900000000000002aa00000000000000fb336e9c1c",
    x"030b00000000000002aafffffffffffff50003e8461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7a71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a9c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fb71c",
    x"070a00000000000002aafffffffffffff8ef35f6ce1c",
    x"080200000000000002aafffffffffffff6f669e1741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfeb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea5f1c",
    x"020900000000000002aa00000000000000fb336e971c",
    x"030b00000000000002aafffffffffffff50003e8471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a991c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fb01c",
    x"070a00000000000002aafffffffffffff8ef35f6cb1c",
    x"080200000000000002aafffffffffffff6f669e1711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfe71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea601c",
    x"020900000000000002aa00000000000000fb336e911c",
    x"030b00000000000002aafffffffffffff50003e8481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a951c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1faa1c",
    x"070a00000000000002aafffffffffffff8ef35f6c71c",
    x"080200000000000002aafffffffffffff6f669e16f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfe31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea621c",
    x"020900000000000002aa00000000000000fb336e8c1c",
    x"030b00000000000002aafffffffffffff50003e8491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc79f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1fa41c",
    x"070a00000000000002aafffffffffffff8ef35f6c31c",
    x"080200000000000002aafffffffffffff6f669e16c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfde1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea631c",
    x"020900000000000002aa00000000000000fb336e861c",
    x"030b00000000000002aafffffffffffff50003e84a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc79d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a8e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1f9e1c",
    x"070a00000000000002aafffffffffffff8ef35f6c01c",
    x"080200000000000002aafffffffffffff6f669e16a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfda1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea641c",
    x"020900000000000002aa00000000000000fb336e801c",
    x"030b00000000000002aafffffffffffff50003e84b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc79b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a8a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1f981c",
    x"070a00000000000002aafffffffffffff8ef35f6bc1c",
    x"080200000000000002aafffffffffffff6f669e1681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfd61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea651c",
    x"020900000000000002aa00000000000000fb336e7b1c",
    x"030b00000000000002aafffffffffffff50003e84c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1f921c",
    x"070a00000000000002aafffffffffffff8ef35f6b81c",
    x"080200000000000002aafffffffffffff6f669e1651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cfd21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea661c",
    x"020900000000000002aa00000000000000fb336e751c",
    x"030b00000000000002aafffffffffffff50003e84d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a831c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1f8b1c",
    x"070a00000000000002aafffffffffffff8ef35f6b51c",
    x"080200000000000002aafffffffffffff6f669e1631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cfce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea671c",
    x"0209000000000000031f00000000000000fb336e6f1c",
    x"030b000000000000031ffffffffffffff50003e84e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc7931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3a7f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1f851c",
    x"070a000000000000031ffffffffffffff8ef35f6b11c",
    x"0802000000000000031ffffffffffffff6f669e1601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cfca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea681c",
    x"020900000000000000ae00000000000000fb336e6a1c",
    x"030b00000000000000aefffffffffffff50003e84f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc7911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3a7c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1f7f1c",
    x"070a00000000000000aefffffffffffff8ef35f6ad1c",
    x"080200000000000000aefffffffffffff6f669e15e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cfc51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea691c",
    x"020900000000000001a400000000000000fb336e641c",
    x"030b00000000000001a4fffffffffffff50003e8501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc78e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3a781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1f791c",
    x"070a00000000000001a4fffffffffffff8ef35f6aa1c",
    x"080200000000000001a4fffffffffffff6f669e15c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266cfc11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbea6b1c",
    x"020900000000000001aa00000000000000fb336e5f1c",
    x"030b00000000000001aafffffffffffff50003e8511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc78c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f3a741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd1f731c",
    x"070a00000000000001aafffffffffffff8ef35f6a61c",
    x"080200000000000001aafffffffffffff6f669e1591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cfbd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbea6c1c",
    x"0209000000000000029500000000000000fb336e591c",
    x"030b0000000000000295fffffffffffff50003e8521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc7891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3a711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1f6d1c",
    x"070a0000000000000295fffffffffffff8ef35f6a21c",
    x"08020000000000000295fffffffffffff6f669e1571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266cfb91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbea6d1c",
    x"0209000000000000015a00000000000000fb336e531c",
    x"030b000000000000015afffffffffffff50003e8521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc7871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3a6d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd1f661c",
    x"070a000000000000015afffffffffffff8ef35f69f1c",
    x"0802000000000000015afffffffffffff6f669e1541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cfb51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbea6e1c",
    x"0209000000000000029500000000000000fb336e4e1c",
    x"030b0000000000000295fffffffffffff50003e8531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc7841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3a691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1f601c",
    x"070a0000000000000295fffffffffffff8ef35f69b1c",
    x"08020000000000000295fffffffffffff6f669e1521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266cfb11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbea6f1c",
    x"0209000000000000015600000000000000fb336e481c",
    x"030b00000000000002aafffffffffffff50003e8541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc7821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd1f5a1c",
    x"070a00000000000002aafffffffffffff8ef35f6971c",
    x"08020000000000000156fffffffffffff6f669e1501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266cfac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea701c",
    x"0209000000000000016500000000000000fb336e431c",
    x"030b000000000000019afffffffffffff50003e8551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc77f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a90000000000000b072f3a621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd1f541c",
    x"070a00000000000001aafffffffffffff8ef35f6941c",
    x"08020000000000000156fffffffffffff6f669e14d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cfa81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbea711c",
    x"020900000000000002a500000000000000fb336e3d1c",
    x"030b000000000000019afffffffffffff50003e8561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc77d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3a5e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd1f4e1c",
    x"070a0000000000000165fffffffffffff8ef35f6901c",
    x"08020000000000000265fffffffffffff6f669e14b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266cfa41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbea721c",
    x"0209000000000000026600000000000000fb336e371c",
    x"030b0000000000000299fffffffffffff50003e8571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc77b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f3a5b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd1f481c",
    x"070a0000000000000256fffffffffffff8ef35f68c1c",
    x"08020000000000000195fffffffffffff6f669e1481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266cfa01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbea741c",
    x"0209000000000000029900000000000000fb336e321c",
    x"030b0000000000000259fffffffffffff50003e8581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc7781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f3a571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd1f411c",
    x"070a0000000000000266fffffffffffff8ef35f6891c",
    x"080200000000000001a5fffffffffffff6f669e1461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266cf9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea751c",
    x"020900000000000002aa00000000000000fb336e2c1c",
    x"030b00000000000002a5fffffffffffff50003e8591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc7761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3a531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd1f3b1c",
    x"070a0000000000000295fffffffffffff8ef35f6851c",
    x"080200000000000001a5fffffffffffff6f669e1441c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266cf971c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbea761c",
    x"020900000000000002a500000000000000fb336e271c",
    x"030b000000000000016afffffffffffff50003e85a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc7731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f3a501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd1f351c",
    x"070a0000000000000255fffffffffffff8ef35f6811c",
    x"08020000000000000169fffffffffffff6f669e1411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266cf931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbea771c",
    x"0209000000000000025600000000000000fb336e211c",
    x"030b0000000000000166fffffffffffff50003e85b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc7711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f3a4c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd1f2f1c",
    x"070a000000000000029afffffffffffff8ef35f67e1c",
    x"08020000000000000295fffffffffffff6f669e13f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000269ffffffffffffff0266cf8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbea781c",
    x"0209000000000000015500000000000000fb336e1b1c",
    x"030b0000000000000296fffffffffffff50003e85c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc76e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3a491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd1f291c",
    x"070a0000000000000156fffffffffffff8ef35f67a1c",
    x"08020000000000000266fffffffffffff6f669e13c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266cf8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbea791c",
    x"0209000000000000016500000000000000fb336e161c",
    x"030b0000000000000265fffffffffffff50003e85d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc76c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3a451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002650000000000000004cd1f231c",
    x"070a0000000000000295fffffffffffff8ef35f6761c",
    x"0802000000000000029afffffffffffff6f669e13a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266cf871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a90000000000000b0bfbea7a1c",
    x"0209000000000000015900000000000000fb336e101c",
    x"030b00000000000002a5fffffffffffff50003e85e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc7691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3a411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002990000000000000004cd1f1c1c",
    x"070a00000000000001a5fffffffffffff8ef35f6731c",
    x"080200000000000001a5fffffffffffff6f669e1381c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266cf831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002690000000000000b0bfbea7b1c",
    x"0209000000000000015500000000000000fb336e0b1c",
    x"030b000000000000019afffffffffffff50003e85f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc7671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f3a3e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002650000000000000004cd1f161c",
    x"070a00000000000002a6fffffffffffff8ef35f66f1c",
    x"08020000000000000256fffffffffffff6f669e1351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266cf7e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea7d1c",
    x"0209000000000000015a00000000000000fb336e051c",
    x"030b00000000000002a5fffffffffffff50003e8601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc7641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3a3a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1f101c",
    x"070a00000000000002a5fffffffffffff8ef35f66b1c",
    x"08020000000000000169fffffffffffff6f669e1331c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cf7a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea7e1c",
    x"0209000000000000031f00000000000000fb336dff1c",
    x"030b000000000000031ffffffffffffff50003e8611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc7621c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f3a361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1f0a1c",
    x"070a000000000000031ffffffffffffff8ef35f6681c",
    x"0802000000000000031ffffffffffffff6f669e1301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cf761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea7f1c",
    x"020900000000000000ae00000000000000fb336dfa1c",
    x"030b00000000000000aefffffffffffff50003e8621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc75f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f3a331c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1f041c",
    x"070a00000000000000aefffffffffffff8ef35f6641c",
    x"080200000000000000aefffffffffffff6f669e12e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cf721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea801c",
    x"020900000000000001a400000000000000fb336df41c",
    x"030b00000000000001a4fffffffffffff50003e8621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc75d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f3a2f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1efe1c",
    x"070a00000000000001a4fffffffffffff8ef35f6601c",
    x"080200000000000001a4fffffffffffff6f669e12c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266cf6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbea811c",
    x"0209000000000000016a00000000000000fb336dee1c",
    x"030b000000000000016afffffffffffff50003e8631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc75b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f3a2b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd1ef71c",
    x"070a000000000000016afffffffffffff8ef35f65c1c",
    x"0802000000000000016afffffffffffff6f669e1291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cf6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea821c",
    x"0209000000000000015500000000000000fb336de91c",
    x"030b0000000000000155fffffffffffff50003e8641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc7581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f3a281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1ef11c",
    x"070a0000000000000155fffffffffffff8ef35f6591c",
    x"08020000000000000155fffffffffffff6f669e1271c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266cf651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbea831c",
    x"0209000000000000019500000000000000fb336de31c",
    x"030b0000000000000195fffffffffffff50003e8651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dc7561c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f3a241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1eeb1c",
    x"070a0000000000000195fffffffffffff8ef35f6551c",
    x"080200000000000002a5fffffffffffff6f669e1241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cf611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea841c",
    x"020900000000000002aa00000000000000fb336dde1c",
    x"030b00000000000002aafffffffffffff50003e8661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1ee51c",
    x"070a00000000000002aafffffffffffff8ef35f6511c",
    x"08020000000000000155fffffffffffff6f669e1221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266cf5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbea861c",
    x"0209000000000000029600000000000000fb336dd81c",
    x"030b00000000000001aafffffffffffff50003e8671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc7511c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f3a1d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd1edf1c",
    x"070a0000000000000256fffffffffffff8ef35f64e1c",
    x"08020000000000000155fffffffffffff6f669e1201c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266cf591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbea871c",
    x"0209000000000000026500000000000000fb336dd21c",
    x"030b00000000000002a9fffffffffffff50003e8681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc74e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3a191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd1ed91c",
    x"070a000000000000029afffffffffffff8ef35f64a1c",
    x"08020000000000000159fffffffffffff6f669e11d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266cf551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbea881c",
    x"0209000000000000029600000000000000fb336dcd1c",
    x"030b000000000000016afffffffffffff50003e8691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc74c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f3a161c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd1ed21c",
    x"070a0000000000000159fffffffffffff8ef35f6461c",
    x"0802000000000000015afffffffffffff6f669e11b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266cf511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea891c",
    x"0209000000000000016900000000000000fb336dc71c",
    x"030b0000000000000295fffffffffffff50003e86a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc7491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f3a121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd1ecc1c",
    x"070a0000000000000196fffffffffffff8ef35f6431c",
    x"08020000000000000299fffffffffffff6f669e1181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266cf4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbea8a1c",
    x"020900000000000002a500000000000000fb336dc21c",
    x"030b0000000000000156fffffffffffff50003e86b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc7471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f3a0e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd1ec61c",
    x"070a00000000000002a6fffffffffffff8ef35f63f1c",
    x"080200000000000001a5fffffffffffff6f669e1161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266cf481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbea8b1c",
    x"0209000000000000025500000000000000fb336dbc1c",
    x"030b000000000000016afffffffffffff50003e86c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc7441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f3a0b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1ec01c",
    x"070a0000000000000295fffffffffffff8ef35f63b1c",
    x"0802000000000000026afffffffffffff6f669e1141c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cf441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbea8c1c",
    x"0209000000000000029a00000000000000fb336db61c",
    x"030b0000000000000269fffffffffffff50003e86d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc7421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f3a071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1eba1c",
    x"070a0000000000000196fffffffffffff8ef35f6381c",
    x"08020000000000000165fffffffffffff6f669e1111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cf401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbea8d1c",
    x"020900000000000001a600000000000000fb336db11c",
    x"030b000000000000019afffffffffffff50003e86e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc73f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f3a031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd1eb41c",
    x"070a000000000000026afffffffffffff8ef35f6341c",
    x"0802000000000000019afffffffffffff6f669e10f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266cf3c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbea8e1c",
    x"0209000000000000025a00000000000000fb336dab1c",
    x"030b00000000000002a9fffffffffffff50003e86f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc73d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f3a001c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd1ead1c",
    x"070a00000000000002a6fffffffffffff8ef35f6301c",
    x"08020000000000000295fffffffffffff6f669e10c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266cf371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbea901c",
    x"0209000000000000029600000000000000fb336da61c",
    x"030b000000000000025afffffffffffff50003e8701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc73a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f39fc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd1ea71c",
    x"070a000000000000019afffffffffffff8ef35f62d1c",
    x"0802000000000000029afffffffffffff6f669e10a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266cf331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbea911c",
    x"0209000000000000019900000000000000fb336da01c",
    x"030b0000000000000156fffffffffffff50003e8711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc7381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f39f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd1ea11c",
    x"070a0000000000000166fffffffffffff8ef35f6291c",
    x"080200000000000001a9fffffffffffff6f669e1081c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266cf2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbea921c",
    x"0209000000000000015600000000000000fb336d9a1c",
    x"030b0000000000000169fffffffffffff50003e8711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc7361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f39f51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd1e9b1c",
    x"070a0000000000000159fffffffffffff8ef35f6251c",
    x"08020000000000000255fffffffffffff6f669e1051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266cf2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbea931c",
    x"0209000000000000029a00000000000000fb336d951c",
    x"030b00000000000002a9fffffffffffff50003e8721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc7331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39f11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd1e951c",
    x"070a0000000000000159fffffffffffff8ef35f6221c",
    x"08020000000000000299fffffffffffff6f669e1031c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cf271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbea941c",
    x"0209000000000000031f00000000000000fb336d8f1c",
    x"030b000000000000031ffffffffffffff50003e8731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc7311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f39ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1e8f1c",
    x"070a000000000000031ffffffffffffff8ef35f61e1c",
    x"0802000000000000031ffffffffffffff6f669e1001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cf231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbea951c",
    x"020900000000000000ae00000000000000fb336d891c",
    x"030b00000000000000aefffffffffffff50003e8741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc72e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f39ea1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1e881c",
    x"070a00000000000000aefffffffffffff8ef35f61a1c",
    x"080200000000000000aefffffffffffff6f669e0fe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cf1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbea961c",
    x"020900000000000001a400000000000000fb336d841c",
    x"030b00000000000001a4fffffffffffff50003e8751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc72c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f39e61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1e821c",
    x"070a00000000000001a4fffffffffffff8ef35f6171c",
    x"080200000000000001a4fffffffffffff6f669e0fc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266cf1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbea971c",
    x"0209000000000000026a00000000000000fb336d7e1c",
    x"030b000000000000026afffffffffffff50003e8761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc7291c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f39e31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026a0000000000000004cd1e7c1c",
    x"070a000000000000026afffffffffffff8ef35f6131c",
    x"0802000000000000026afffffffffffff6f669e0f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cf161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea991c",
    x"020900000000000002aa00000000000000fb336d791c",
    x"030b00000000000002aafffffffffffff50003e8771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f39df1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd1e761c",
    x"070a0000000000000156fffffffffffff8ef35f60f1c",
    x"080200000000000002aafffffffffffff6f669e0f71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cf121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbea9a1c",
    x"020900000000000002aa00000000000000fb336d731c",
    x"030b00000000000002aafffffffffffff50003e8781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39db1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1e701c",
    x"070a0000000000000255fffffffffffff8ef35f60c1c",
    x"080200000000000002aafffffffffffff6f669e0f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266cf0e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbea9b1c",
    x"020900000000000002a900000000000000fb336d6d1c",
    x"030b00000000000002aafffffffffffff50003e8791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a9fffffffffffff4099dc7221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f39d81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd1e6a1c",
    x"070a0000000000000155fffffffffffff8ef35f6081c",
    x"080200000000000002aafffffffffffff6f669e0f21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cf0a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a90000000000000b0bfbea9c1c",
    x"020900000000000001aa00000000000000fb336d681c",
    x"030b000000000000026afffffffffffff50003e87a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc71f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f39d41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd1e631c",
    x"070a0000000000000195fffffffffffff8ef35f6041c",
    x"0802000000000000026afffffffffffff6f669e0f01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266cf051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbea9d1c",
    x"0209000000000000029a00000000000000fb336d621c",
    x"030b0000000000000156fffffffffffff50003e87b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc71d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39d01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd1e5d1c",
    x"070a00000000000001a9fffffffffffff8ef35f6011c",
    x"08020000000000000166fffffffffffff6f669e0ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266cf011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbea9e1c",
    x"0209000000000000026600000000000000fb336d5d1c",
    x"030b000000000000026afffffffffffff50003e87c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc71a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f39cd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd1e571c",
    x"070a0000000000000199fffffffffffff8ef35f5fd1c",
    x"08020000000000000159fffffffffffff6f669e0eb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000299ffffffffffffff0266cefd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbea9f1c",
    x"0209000000000000029a00000000000000fb336d571c",
    x"030b0000000000000299fffffffffffff50003e87d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc7181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f39c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd1e511c",
    x"070a00000000000002a9fffffffffffff8ef35f5f91c",
    x"080200000000000001a5fffffffffffff6f669e0e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266cef91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbeaa01c",
    x"0209000000000000026a00000000000000fb336d511c",
    x"030b000000000000019afffffffffffff50003e87e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc7151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f39c51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd1e4b1c",
    x"070a00000000000001a5fffffffffffff8ef35f5f61c",
    x"08020000000000000295fffffffffffff6f669e0e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cef51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbeaa21c",
    x"0209000000000000019500000000000000fb336d4c1c",
    x"030b0000000000000155fffffffffffff50003e87f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc7131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f39c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd1e451c",
    x"070a000000000000026afffffffffffff8ef35f5f21c",
    x"0802000000000000026afffffffffffff6f669e0e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266cef01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbeaa31c",
    x"020900000000000001a900000000000000fb336d461c",
    x"030b000000000000015afffffffffffff50003e8801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dc7111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f39be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd1e3e1c",
    x"070a000000000000015afffffffffffff8ef35f5ee1c",
    x"0802000000000000016afffffffffffff6f669e0e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266ceec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbeaa41c",
    x"0209000000000000025600000000000000fb336d411c",
    x"030b00000000000002aafffffffffffff50003e8801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc70e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f39ba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd1e381c",
    x"070a00000000000001a9fffffffffffff8ef35f5eb1c",
    x"08020000000000000266fffffffffffff6f669e0df1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266cee81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbeaa51c",
    x"0209000000000000016a00000000000000fb336d3b1c",
    x"030b0000000000000166fffffffffffff50003e8811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc70c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f39b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd1e321c",
    x"070a0000000000000199fffffffffffff8ef35f5e71c",
    x"08020000000000000299fffffffffffff6f669e0dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266cee41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbeaa61c",
    x"0209000000000000029600000000000000fb336d351c",
    x"030b0000000000000295fffffffffffff50003e8821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc7091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f39b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd1e2c1c",
    x"070a00000000000001a9fffffffffffff8ef35f5e31c",
    x"08020000000000000266fffffffffffff6f669e0da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266cee01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbeaa71c",
    x"0209000000000000019500000000000000fb336d301c",
    x"030b0000000000000295fffffffffffff50003e8831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000259fffffffffffff4099dc7071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f39b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd1e261c",
    x"070a000000000000025afffffffffffff8ef35f5e01c",
    x"08020000000000000199fffffffffffff6f669e0d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cedc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbeaa81c",
    x"0209000000000000015600000000000000fb336d2a1c",
    x"030b0000000000000295fffffffffffff50003e8841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc7041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f39ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001990000000000000004cd1e201c",
    x"070a0000000000000199fffffffffffff8ef35f5dc1c",
    x"08020000000000000269fffffffffffff6f669e0d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266ced71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbeaa91c",
    x"020900000000000002a600000000000000fb336d251c",
    x"030b000000000000015afffffffffffff50003e8851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc7021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f39a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002990000000000000004cd1e191c",
    x"070a0000000000000295fffffffffffff8ef35f5d81c",
    x"080200000000000002a5fffffffffffff6f669e0d31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266ced31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeaab1c",
    x"0209000000000000031f00000000000000fb336d1f1c",
    x"030b000000000000031ffffffffffffff50003e8861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc6ff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f39a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1e131c",
    x"070a000000000000031ffffffffffffff8ef35f5d51c",
    x"0802000000000000031ffffffffffffff6f669e0d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cecf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeaac1c",
    x"020900000000000000ae00000000000000fb336d191c",
    x"030b00000000000000aefffffffffffff50003e8871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc6fd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f39a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1e0d1c",
    x"070a00000000000000aefffffffffffff8ef35f5d11c",
    x"080200000000000000aefffffffffffff6f669e0ce1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cecb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeaad1c",
    x"020900000000000001a400000000000000fb336d141c",
    x"030b00000000000001a4fffffffffffff50003e8881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc6fa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f399d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1e071c",
    x"070a00000000000001a4fffffffffffff8ef35f5cd1c",
    x"080200000000000001a4fffffffffffff6f669e0cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266cec71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbeaae1c",
    x"0209000000000000015a00000000000000fb336d0e1c",
    x"030b000000000000015afffffffffffff50003e8891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc6f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f399a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd1e011c",
    x"070a000000000000015afffffffffffff8ef35f5ca1c",
    x"0802000000000000015afffffffffffff6f669e0c91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cec31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeaaf1c",
    x"020900000000000001aa00000000000000fb336d081c",
    x"030b0000000000000255fffffffffffff50003e88a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6f51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1dfb1c",
    x"070a0000000000000155fffffffffffff8ef35f5c61c",
    x"08020000000000000155fffffffffffff6f669e0c71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266cebe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbeab01c",
    x"0209000000000000016900000000000000fb336d031c",
    x"030b0000000000000269fffffffffffff50003e88b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc6f31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f39921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd1df41c",
    x"070a00000000000002a6fffffffffffff8ef35f5c21c",
    x"080200000000000001a5fffffffffffff6f669e0c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266ceba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbeab11c",
    x"020900000000000001a600000000000000fb336cfd1c",
    x"030b0000000000000296fffffffffffff50003e88c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc6f01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f398f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd1dee1c",
    x"070a000000000000029afffffffffffff8ef35f5bf1c",
    x"08020000000000000196fffffffffffff6f669e0c21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266ceb61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbeab21c",
    x"0209000000000000026900000000000000fb336cf81c",
    x"030b0000000000000255fffffffffffff50003e88d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc6ee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f398b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001990000000000000004cd1de81c",
    x"070a0000000000000265fffffffffffff8ef35f5bb1c",
    x"08020000000000000256fffffffffffff6f669e0bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ceb21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbeab41c",
    x"0209000000000000015600000000000000fb336cf21c",
    x"030b0000000000000155fffffffffffff50003e88e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f39871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd1de21c",
    x"070a00000000000002aafffffffffffff8ef35f5b71c",
    x"08020000000000000155fffffffffffff6f669e0bd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266ceae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbeab51c",
    x"0209000000000000026500000000000000fb336cec1c",
    x"030b0000000000000265fffffffffffff50003e88e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc6e91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f39841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002650000000000000004cd1ddc1c",
    x"070a000000000000019afffffffffffff8ef35f5b41c",
    x"08020000000000000265fffffffffffff6f669e0bb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ceaa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeab61c",
    x"0209000000000000015500000000000000fb336ce71c",
    x"030b0000000000000155fffffffffffff50003e88f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6e71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1dd61c",
    x"070a00000000000002aafffffffffffff8ef35f5b01c",
    x"08020000000000000155fffffffffffff6f669e0b81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cea51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeab71c",
    x"0209000000000000015500000000000000fb336ce11c",
    x"030b0000000000000155fffffffffffff50003e8901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f397d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1dcf1c",
    x"070a00000000000002aafffffffffffff8ef35f5ac1c",
    x"08020000000000000155fffffffffffff6f669e0b61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cea11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeab81c",
    x"0209000000000000015500000000000000fb336cdc1c",
    x"030b0000000000000155fffffffffffff50003e8911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6e21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1dc91c",
    x"070a00000000000002aafffffffffffff8ef35f5a91c",
    x"08020000000000000155fffffffffffff6f669e0b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266ce9d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbeab91c",
    x"0209000000000000025900000000000000fb336cd61c",
    x"030b0000000000000259fffffffffffff50003e8921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc6df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f39751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002590000000000000004cd1dc31c",
    x"070a00000000000001a6fffffffffffff8ef35f5a51c",
    x"08020000000000000259fffffffffffff6f669e0b11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeaba1c",
    x"0209000000000000015500000000000000fb336cd01c",
    x"030b0000000000000155fffffffffffff50003e8931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6dd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1dbd1c",
    x"070a00000000000002aafffffffffffff8ef35f5a11c",
    x"08020000000000000155fffffffffffff6f669e0af1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeabb1c",
    x"0209000000000000015500000000000000fb336ccb1c",
    x"030b0000000000000155fffffffffffff50003e8941c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f396e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1db71c",
    x"070a00000000000002aafffffffffffff8ef35f59e1c",
    x"08020000000000000155fffffffffffff6f669e0ac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266ce911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbeabd1c",
    x"0209000000000000015900000000000000fb336cc51c",
    x"030b0000000000000159fffffffffffff50003e8951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc6d81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f396a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd1db11c",
    x"070a00000000000002a6fffffffffffff8ef35f59a1c",
    x"08020000000000000159fffffffffffff6f669e0aa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266ce8c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbeabe1c",
    x"0209000000000000016a00000000000000fb336cc01c",
    x"030b0000000000000155fffffffffffff50003e8961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc6d51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f39671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1daa1c",
    x"070a0000000000000265fffffffffffff8ef35f5961c",
    x"0802000000000000015afffffffffffff6f669e0a71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266ce881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbeabf1c",
    x"0209000000000000025500000000000000fb336cba1c",
    x"030b0000000000000255fffffffffffff50003e8971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dc6d31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f39631c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd1da41c",
    x"070a000000000000015afffffffffffff8ef35f5931c",
    x"08020000000000000295fffffffffffff6f669e0a51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266ce841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbeac01c",
    x"020900000000000002a600000000000000fb336cb41c",
    x"030b00000000000002a6fffffffffffff50003e8981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc6d01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f395f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd1d9e1c",
    x"070a0000000000000159fffffffffffff8ef35f58f1c",
    x"080200000000000002a6fffffffffffff6f669e0a31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266ce801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeac11c",
    x"0209000000000000031f00000000000000fb336caf1c",
    x"030b000000000000031ffffffffffffff50003e8991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc6ce1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f395c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1d981c",
    x"070a000000000000031ffffffffffffff8ef35f58b1c",
    x"0802000000000000031ffffffffffffff6f669e0a01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266ce7c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeac21c",
    x"020900000000000000ae00000000000000fb336ca91c",
    x"030b00000000000000aefffffffffffff50003e89a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc6cb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f39581c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1d921c",
    x"070a00000000000000aefffffffffffff8ef35f5871c",
    x"080200000000000000aefffffffffffff6f669e09e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ce771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeac31c",
    x"020900000000000001a400000000000000fb336ca31c",
    x"030b00000000000001a4fffffffffffff50003e89b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc6c91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f39551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1d8c1c",
    x"070a00000000000001a4fffffffffffff8ef35f5841c",
    x"080200000000000001a4fffffffffffff6f669e09b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266ce731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbeac41c",
    x"0209000000000000025a00000000000000fb336c9e1c",
    x"030b000000000000025afffffffffffff50003e89c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc6c61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f39511c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd1d851c",
    x"070a000000000000025afffffffffffff8ef35f5801c",
    x"0802000000000000025afffffffffffff6f669e0991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce6f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeac61c",
    x"020900000000000002aa00000000000000fb336c981c",
    x"030b00000000000002aafffffffffffff50003e89c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6c41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f394d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d7f1c",
    x"070a00000000000002aafffffffffffff8ef35f57c1c",
    x"080200000000000002aafffffffffffff6f669e0971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266ce6b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbeac71c",
    x"0209000000000000029a00000000000000fb336c931c",
    x"030b000000000000029afffffffffffff50003e89d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc6c11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f394a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd1d791c",
    x"070a000000000000029afffffffffffff8ef35f5791c",
    x"0802000000000000029afffffffffffff6f669e0941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeac81c",
    x"020900000000000002aa00000000000000fb336c8d1c",
    x"030b00000000000002aafffffffffffff50003e89e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6bf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39461c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d731c",
    x"070a00000000000002aafffffffffffff8ef35f5751c",
    x"080200000000000002aafffffffffffff6f669e0921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeac91c",
    x"020900000000000002aa00000000000000fb336c871c",
    x"030b00000000000002aafffffffffffff50003e89f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d6d1c",
    x"070a00000000000002aafffffffffffff8ef35f5711c",
    x"080200000000000002aafffffffffffff6f669e08f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce5e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeaca1c",
    x"020900000000000002aa00000000000000fb336c821c",
    x"030b00000000000002aafffffffffffff50003e8a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6ba1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f393f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d671c",
    x"070a00000000000002aafffffffffffff8ef35f56e1c",
    x"080200000000000002aafffffffffffff6f669e08d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce5a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeacb1c",
    x"020900000000000002aa00000000000000fb336c7c1c",
    x"030b00000000000002aafffffffffffff50003e8a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f393b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d601c",
    x"070a00000000000002aafffffffffffff8ef35f56a1c",
    x"080200000000000002aafffffffffffff6f669e08b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeacc1c",
    x"020900000000000002aa00000000000000fb336c771c",
    x"030b00000000000002aafffffffffffff50003e8a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6b51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d5a1c",
    x"070a00000000000002aafffffffffffff8ef35f5661c",
    x"080200000000000002aafffffffffffff6f669e0881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeacd1c",
    x"020900000000000002aa00000000000000fb336c711c",
    x"030b00000000000002aafffffffffffff50003e8a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d541c",
    x"070a00000000000002aafffffffffffff8ef35f5631c",
    x"080200000000000002aafffffffffffff6f669e0861c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce4e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeacf1c",
    x"020900000000000002aa00000000000000fb336c6b1c",
    x"030b00000000000002aafffffffffffff50003e8a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6b01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39301c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d4e1c",
    x"070a00000000000002aafffffffffffff8ef35f55f1c",
    x"080200000000000002aafffffffffffff6f669e0831c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266ce4a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbead01c",
    x"0209000000000000016600000000000000fb336c661c",
    x"030b0000000000000166fffffffffffff50003e8a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc6ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f392d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd1d481c",
    x"070a0000000000000166fffffffffffff8ef35f55b1c",
    x"08020000000000000166fffffffffffff6f669e0811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce451c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbead11c",
    x"0209000000000000015500000000000000fb336c601c",
    x"030b0000000000000155fffffffffffff50003e8a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6ab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1d411c",
    x"070a0000000000000155fffffffffffff8ef35f5581c",
    x"08020000000000000155fffffffffffff6f669e07e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce411c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbead21c",
    x"0209000000000000015500000000000000fb336c5b1c",
    x"030b0000000000000155fffffffffffff50003e8a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39251c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1d3b1c",
    x"070a0000000000000155fffffffffffff8ef35f5541c",
    x"08020000000000000155fffffffffffff6f669e07c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce3d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbead31c",
    x"0209000000000000015500000000000000fb336c551c",
    x"030b0000000000000155fffffffffffff50003e8a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6a61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39221c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1d351c",
    x"070a0000000000000155fffffffffffff8ef35f5501c",
    x"08020000000000000155fffffffffffff6f669e07a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbead41c",
    x"0209000000000000015500000000000000fb336c4f1c",
    x"030b0000000000000155fffffffffffff50003e8a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f391e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1d2f1c",
    x"070a0000000000000155fffffffffffff8ef35f54d1c",
    x"08020000000000000155fffffffffffff6f669e0771c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbead51c",
    x"0209000000000000015500000000000000fb336c4a1c",
    x"030b0000000000000155fffffffffffff50003e8aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6a11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f391a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1d291c",
    x"070a0000000000000155fffffffffffff8ef35f5491c",
    x"08020000000000000155fffffffffffff6f669e0751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266ce311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbead61c",
    x"0209000000000000015900000000000000fb336c441c",
    x"030b0000000000000159fffffffffffff50003e8aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc69f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f39171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd1d231c",
    x"070a0000000000000159fffffffffffff8ef35f5451c",
    x"08020000000000000159fffffffffffff6f669e0721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266ce2c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbead71c",
    x"0209000000000000031f00000000000000fb336c3f1c",
    x"030b000000000000031ffffffffffffff50003e8ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc69c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f39131c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1d1c1c",
    x"070a000000000000031ffffffffffffff8ef35f5421c",
    x"0802000000000000031ffffffffffffff6f669e0701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266ce281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbead91c",
    x"020900000000000000ae00000000000000fb336c391c",
    x"030b00000000000000aefffffffffffff50003e8ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc69a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f390f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1d161c",
    x"070a00000000000000aefffffffffffff8ef35f53e1c",
    x"080200000000000000aefffffffffffff6f669e06e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ce241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeada1c",
    x"020900000000000001a400000000000000fb336c331c",
    x"030b00000000000001a4fffffffffffff50003e8ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc6971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f390c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1d101c",
    x"070a00000000000001a4fffffffffffff8ef35f53a1c",
    x"080200000000000001a4fffffffffffff6f669e06b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266ce201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbeadb1c",
    x"0209000000000000029a00000000000000fb336c2e1c",
    x"030b000000000000029afffffffffffff50003e8ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc6951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f39081c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd1d0a1c",
    x"070a000000000000029afffffffffffff8ef35f5371c",
    x"0802000000000000029afffffffffffff6f669e0691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ce1c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeadc1c",
    x"020900000000000002aa00000000000000fb336c281c",
    x"030b00000000000002aafffffffffffff50003e8af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc6921c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f39051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1d041c",
    x"070a00000000000002aafffffffffffff8ef35f5331c",
    x"080200000000000002aafffffffffffff6f669e0661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeadd1c",
    x"0209000000000000015500000000000000fb336c221c",
    x"030b0000000000000155fffffffffffff50003e8b01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f39011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cfe1c",
    x"070a0000000000000155fffffffffffff8ef35f52f1c",
    x"08020000000000000155fffffffffffff6f669e0641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce131c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeade1c",
    x"0209000000000000015500000000000000fb336c1d1c",
    x"030b0000000000000155fffffffffffff50003e8b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc68e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38fd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cf71c",
    x"070a0000000000000155fffffffffffff8ef35f52c1c",
    x"08020000000000000155fffffffffffff6f669e0621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce0f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeadf1c",
    x"0209000000000000015500000000000000fb336c171c",
    x"030b0000000000000155fffffffffffff50003e8b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc68b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38fa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cf11c",
    x"070a0000000000000155fffffffffffff8ef35f5281c",
    x"08020000000000000155fffffffffffff6f669e05f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce0b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae01c",
    x"0209000000000000015500000000000000fb336c121c",
    x"030b0000000000000155fffffffffffff50003e8b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38f61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1ceb1c",
    x"070a0000000000000155fffffffffffff8ef35f5241c",
    x"08020000000000000155fffffffffffff6f669e05d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae21c",
    x"0209000000000000015500000000000000fb336c0c1c",
    x"030b0000000000000155fffffffffffff50003e8b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38f21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1ce51c",
    x"070a0000000000000155fffffffffffff8ef35f5211c",
    x"08020000000000000155fffffffffffff6f669e05a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ce031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae31c",
    x"0209000000000000015500000000000000fb336c061c",
    x"030b0000000000000155fffffffffffff50003e8b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38ef1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cdf1c",
    x"070a0000000000000155fffffffffffff8ef35f51d1c",
    x"08020000000000000155fffffffffffff6f669e0581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdfe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae41c",
    x"0209000000000000015500000000000000fb336c011c",
    x"030b0000000000000155fffffffffffff50003e8b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cd91c",
    x"070a0000000000000155fffffffffffff8ef35f5191c",
    x"08020000000000000155fffffffffffff6f669e0561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdfa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae51c",
    x"0209000000000000015500000000000000fb336bfb1c",
    x"030b0000000000000155fffffffffffff50003e8b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc67f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38e71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cd21c",
    x"070a0000000000000155fffffffffffff8ef35f5151c",
    x"08020000000000000155fffffffffffff6f669e0531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdf61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae61c",
    x"0209000000000000015500000000000000fb336bf61c",
    x"030b0000000000000155fffffffffffff50003e8b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc67c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38e41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1ccc1c",
    x"070a0000000000000155fffffffffffff8ef35f5121c",
    x"08020000000000000155fffffffffffff6f669e0511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdf21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae71c",
    x"0209000000000000015500000000000000fb336bf01c",
    x"030b0000000000000155fffffffffffff50003e8b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc67a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38e01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cc61c",
    x"070a0000000000000155fffffffffffff8ef35f50e1c",
    x"08020000000000000155fffffffffffff6f669e04e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae81c",
    x"0209000000000000015500000000000000fb336bea1c",
    x"030b0000000000000155fffffffffffff50003e8b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38dd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cc01c",
    x"070a0000000000000155fffffffffffff8ef35f50a1c",
    x"08020000000000000155fffffffffffff6f669e04c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeae91c",
    x"0209000000000000015500000000000000fb336be51c",
    x"030b0000000000000155fffffffffffff50003e8ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cba1c",
    x"070a0000000000000155fffffffffffff8ef35f5071c",
    x"08020000000000000155fffffffffffff6f669e04a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cde51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaeb1c",
    x"0209000000000000015500000000000000fb336bdf1c",
    x"030b0000000000000155fffffffffffff50003e8bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6721c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38d51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1cb41c",
    x"070a0000000000000155fffffffffffff8ef35f5031c",
    x"08020000000000000155fffffffffffff6f669e0471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cde11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbeaec1c",
    x"0209000000000000029500000000000000fb336bda1c",
    x"030b0000000000000295fffffffffffff50003e8bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc6701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f38d21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1cad1c",
    x"070a0000000000000295fffffffffffff8ef35f4ff1c",
    x"08020000000000000295fffffffffffff6f669e0451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cddd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaed1c",
    x"0209000000000000015500000000000000fb336bd41c",
    x"030b0000000000000155fffffffffffff50003e8bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc66d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1ca71c",
    x"070a0000000000000155fffffffffffff8ef35f4fc1c",
    x"08020000000000000155fffffffffffff6f669e0421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cdd91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeaee1c",
    x"0209000000000000031f00000000000000fb336bce1c",
    x"030b000000000000031ffffffffffffff50003e8be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc66b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f38ca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1ca11c",
    x"070a000000000000031ffffffffffffff8ef35f4f81c",
    x"0802000000000000031ffffffffffffff6f669e0401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cdd51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeaef1c",
    x"020900000000000000ae00000000000000fb336bc91c",
    x"030b00000000000000aefffffffffffff50003e8bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc6681c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f38c71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1c9b1c",
    x"070a00000000000000aefffffffffffff8ef35f4f41c",
    x"080200000000000000aefffffffffffff6f669e03e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cdd11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeaf01c",
    x"020900000000000001a400000000000000fb336bc31c",
    x"030b00000000000001a4fffffffffffff50003e8c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc6661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f38c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1c951c",
    x"070a00000000000001a4fffffffffffff8ef35f4f11c",
    x"080200000000000001a4fffffffffffff6f669e03b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266cdcc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbeaf11c",
    x"0209000000000000019a00000000000000fb336bbd1c",
    x"030b000000000000019afffffffffffff50003e8c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc6631c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f38bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd1c8f1c",
    x"070a000000000000019afffffffffffff8ef35f4ed1c",
    x"0802000000000000019afffffffffffff6f669e0391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdc81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf21c",
    x"0209000000000000015500000000000000fb336bb81c",
    x"030b0000000000000155fffffffffffff50003e8c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38bc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c881c",
    x"070a0000000000000155fffffffffffff8ef35f4e91c",
    x"08020000000000000155fffffffffffff6f669e0361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdc41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf41c",
    x"0209000000000000015500000000000000fb336bb21c",
    x"030b0000000000000155fffffffffffff50003e8c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc65f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38b81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c821c",
    x"070a0000000000000155fffffffffffff8ef35f4e61c",
    x"08020000000000000155fffffffffffff6f669e0341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdc01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf51c",
    x"0209000000000000015500000000000000fb336bad1c",
    x"030b0000000000000155fffffffffffff50003e8c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc65c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38b51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c7c1c",
    x"070a0000000000000155fffffffffffff8ef35f4e21c",
    x"08020000000000000155fffffffffffff6f669e0311c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdbc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf61c",
    x"0209000000000000015500000000000000fb336ba71c",
    x"030b0000000000000155fffffffffffff50003e8c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc65a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38b11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c761c",
    x"070a0000000000000155fffffffffffff8ef35f4de1c",
    x"08020000000000000155fffffffffffff6f669e02f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdb81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf71c",
    x"0209000000000000015500000000000000fb336ba11c",
    x"030b0000000000000155fffffffffffff50003e8c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38ad1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c701c",
    x"070a0000000000000155fffffffffffff8ef35f4db1c",
    x"08020000000000000155fffffffffffff6f669e02d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdb31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf81c",
    x"0209000000000000015500000000000000fb336b9c1c",
    x"030b0000000000000155fffffffffffff50003e8c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38aa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c6a1c",
    x"070a0000000000000155fffffffffffff8ef35f4d71c",
    x"08020000000000000155fffffffffffff6f669e02a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdaf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaf91c",
    x"0209000000000000015500000000000000fb336b961c",
    x"030b0000000000000155fffffffffffff50003e8c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38a61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c631c",
    x"070a0000000000000155fffffffffffff8ef35f4d31c",
    x"08020000000000000155fffffffffffff6f669e0281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cdab1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeafa1c",
    x"0209000000000000015500000000000000fb336b911c",
    x"030b0000000000000155fffffffffffff50003e8c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38a21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c5d1c",
    x"070a0000000000000155fffffffffffff8ef35f4d01c",
    x"08020000000000000155fffffffffffff6f669e0251c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cda71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeafb1c",
    x"0209000000000000015500000000000000fb336b8b1c",
    x"030b0000000000000155fffffffffffff50003e8c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc64d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f389f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c571c",
    x"070a0000000000000155fffffffffffff8ef35f4cc1c",
    x"08020000000000000155fffffffffffff6f669e0231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cda31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeafd1c",
    x"0209000000000000015500000000000000fb336b851c",
    x"030b0000000000000155fffffffffffff50003e8ca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc64b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f389b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c511c",
    x"070a0000000000000155fffffffffffff8ef35f4c81c",
    x"08020000000000000155fffffffffffff6f669e0211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd9e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeafe1c",
    x"0209000000000000015500000000000000fb336b801c",
    x"030b0000000000000155fffffffffffff50003e8cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38971c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c4b1c",
    x"070a0000000000000155fffffffffffff8ef35f4c51c",
    x"08020000000000000155fffffffffffff6f669e01e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd9a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeaff1c",
    x"0209000000000000015500000000000000fb336b7a1c",
    x"030b0000000000000155fffffffffffff50003e8cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c451c",
    x"070a0000000000000155fffffffffffff8ef35f4c11c",
    x"08020000000000000155fffffffffffff6f669e01c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd961c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb001c",
    x"0209000000000000015500000000000000fb336b751c",
    x"030b0000000000000155fffffffffffff50003e8cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38901c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c3e1c",
    x"070a0000000000000155fffffffffffff8ef35f4bd1c",
    x"08020000000000000155fffffffffffff6f669e0191c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd921c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb011c",
    x"0209000000000000015500000000000000fb336b6f1c",
    x"030b0000000000000155fffffffffffff50003e8ce1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f388d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c381c",
    x"070a0000000000000155fffffffffffff8ef35f4b91c",
    x"08020000000000000155fffffffffffff6f669e0171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd8e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb021c",
    x"0209000000000000015500000000000000fb336b691c",
    x"030b0000000000000155fffffffffffff50003e8cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc63e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c321c",
    x"070a0000000000000155fffffffffffff8ef35f4b61c",
    x"08020000000000000155fffffffffffff6f669e0151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd8a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb031c",
    x"0209000000000000015500000000000000fb336b641c",
    x"030b0000000000000155fffffffffffff50003e8d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc63c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38851c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c2c1c",
    x"070a0000000000000155fffffffffffff8ef35f4b21c",
    x"08020000000000000155fffffffffffff6f669e0121c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cd851c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb041c",
    x"0209000000000000031f00000000000000fb336b5e1c",
    x"030b000000000000031ffffffffffffff50003e8d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc6391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f38821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1c261c",
    x"070a000000000000031ffffffffffffff8ef35f4ae1c",
    x"0802000000000000031ffffffffffffff6f669e0101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cd811c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb061c",
    x"020900000000000000ae00000000000000fb336b581c",
    x"030b00000000000000aefffffffffffff50003e8d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc6371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f387e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1c1f1c",
    x"070a00000000000000aefffffffffffff8ef35f4ab1c",
    x"080200000000000000aefffffffffffff6f669e00d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cd7d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb071c",
    x"020900000000000001a400000000000000fb336b531c",
    x"030b00000000000001a4fffffffffffff50003e8d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc6341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f387a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1c191c",
    x"070a00000000000001a4fffffffffffff8ef35f4a71c",
    x"080200000000000001a4fffffffffffff6f669e00b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266cd791c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbeb081c",
    x"0209000000000000015600000000000000fb336b4d1c",
    x"030b0000000000000156fffffffffffff50003e8d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc6321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f38771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd1c131c",
    x"070a0000000000000156fffffffffffff8ef35f4a31c",
    x"08020000000000000156fffffffffffff6f669e0091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cd751c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbeb091c",
    x"0209000000000000029500000000000000fb336b481c",
    x"030b0000000000000295fffffffffffff50003e8d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc62f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f38731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1c0d1c",
    x"070a0000000000000295fffffffffffff8ef35f4a01c",
    x"08020000000000000295fffffffffffff6f669e0061c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266cd711c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbeb0a1c",
    x"0209000000000000016600000000000000fb336b421c",
    x"030b0000000000000166fffffffffffff50003e8d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc62d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f386f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd1c071c",
    x"070a0000000000000166fffffffffffff8ef35f49c1c",
    x"08020000000000000166fffffffffffff6f669e0041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd6c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb0b1c",
    x"0209000000000000015500000000000000fb336b3c1c",
    x"030b0000000000000155fffffffffffff50003e8d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc62b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f386c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1c011c",
    x"070a0000000000000155fffffffffffff8ef35f4981c",
    x"08020000000000000155fffffffffffff6f669e0011c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd681c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb0c1c",
    x"0209000000000000015500000000000000fb336b371c",
    x"030b0000000000000155fffffffffffff50003e8d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bfa1c",
    x"070a0000000000000155fffffffffffff8ef35f4951c",
    x"08020000000000000155fffffffffffff6f669dfff1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd641c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb0e1c",
    x"0209000000000000015500000000000000fb336b311c",
    x"030b0000000000000155fffffffffffff50003e8d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bf41c",
    x"070a0000000000000155fffffffffffff8ef35f4911c",
    x"08020000000000000155fffffffffffff6f669dffd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd601c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb0f1c",
    x"0209000000000000015500000000000000fb336b2c1c",
    x"030b0000000000000155fffffffffffff50003e8d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bee1c",
    x"070a0000000000000155fffffffffffff8ef35f48d1c",
    x"08020000000000000155fffffffffffff6f669dffa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd5c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb101c",
    x"0209000000000000015500000000000000fb336b261c",
    x"030b0000000000000155fffffffffffff50003e8da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f385d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1be81c",
    x"070a0000000000000155fffffffffffff8ef35f48a1c",
    x"08020000000000000155fffffffffffff6f669dff81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd581c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb111c",
    x"0209000000000000015500000000000000fb336b201c",
    x"030b0000000000000155fffffffffffff50003e8db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc61e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f385a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1be21c",
    x"070a0000000000000155fffffffffffff8ef35f4861c",
    x"08020000000000000155fffffffffffff6f669dff51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd531c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb121c",
    x"0209000000000000015500000000000000fb336b1b1c",
    x"030b0000000000000155fffffffffffff50003e8dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc61c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bdc1c",
    x"070a0000000000000155fffffffffffff8ef35f4821c",
    x"08020000000000000155fffffffffffff6f669dff31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd4f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb131c",
    x"0209000000000000015500000000000000fb336b151c",
    x"030b0000000000000155fffffffffffff50003e8dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bd51c",
    x"070a0000000000000155fffffffffffff8ef35f47f1c",
    x"08020000000000000155fffffffffffff6f669dff01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd4b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb141c",
    x"0209000000000000015500000000000000fb336b101c",
    x"030b0000000000000155fffffffffffff50003e8de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f384f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bcf1c",
    x"070a0000000000000155fffffffffffff8ef35f47b1c",
    x"08020000000000000155fffffffffffff6f669dfee1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd471c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb151c",
    x"0209000000000000015500000000000000fb336b0a1c",
    x"030b0000000000000155fffffffffffff50003e8de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f384b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bc91c",
    x"070a0000000000000155fffffffffffff8ef35f4771c",
    x"08020000000000000155fffffffffffff6f669dfec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd431c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb171c",
    x"0209000000000000015500000000000000fb336b041c",
    x"030b0000000000000155fffffffffffff50003e8df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc6121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bc31c",
    x"070a0000000000000155fffffffffffff8ef35f4741c",
    x"08020000000000000155fffffffffffff6f669dfe91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd3f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb181c",
    x"0209000000000000015500000000000000fb336aff1c",
    x"030b0000000000000155fffffffffffff50003e8e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc60f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f38441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bbd1c",
    x"070a0000000000000155fffffffffffff8ef35f4701c",
    x"08020000000000000155fffffffffffff6f669dfe71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cd3a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbeb191c",
    x"0209000000000000029500000000000000fb336af91c",
    x"030b0000000000000295fffffffffffff50003e8e11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc60d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f38401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd1bb71c",
    x"070a0000000000000295fffffffffffff8ef35f46c1c",
    x"08020000000000000295fffffffffffff6f669dfe41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cd361c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb1a1c",
    x"0209000000000000015500000000000000fb336af31c",
    x"030b0000000000000155fffffffffffff50003e8e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc60a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f383d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1bb01c",
    x"070a0000000000000155fffffffffffff8ef35f4681c",
    x"08020000000000000155fffffffffffff6f669dfe21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cd321c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb1b1c",
    x"0209000000000000031f00000000000000fb336aee1c",
    x"030b000000000000031ffffffffffffff50003e8e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc6081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f38391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1baa1c",
    x"070a000000000000031ffffffffffffff8ef35f4651c",
    x"0802000000000000031ffffffffffffff6f669dfe01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cd2e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb1c1c",
    x"020900000000000000ae00000000000000fb336ae81c",
    x"030b00000000000000aefffffffffffff50003e8e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc6051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f38351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1ba41c",
    x"070a00000000000000aefffffffffffff8ef35f4611c",
    x"080200000000000000aefffffffffffff6f669dfdd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cd2a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb1d1c",
    x"020900000000000001a400000000000000fb336ae31c",
    x"030b00000000000001a4fffffffffffff50003e8e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc6031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f38321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1b9e1c",
    x"070a00000000000001a4fffffffffffff8ef35f45d1c",
    x"080200000000000001a4fffffffffffff6f669dfdb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266cd261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbeb1e1c",
    x"0209000000000000025600000000000000fb336add1c",
    x"030b0000000000000256fffffffffffff50003e8e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dc6001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f382e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd1b981c",
    x"070a0000000000000256fffffffffffff8ef35f45a1c",
    x"08020000000000000256fffffffffffff6f669dfd81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb201c",
    x"020900000000000002aa00000000000000fb336ad71c",
    x"030b00000000000002aafffffffffffff50003e8e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5fe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f382a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b921c",
    x"070a00000000000002aafffffffffffff8ef35f4561c",
    x"080200000000000002aafffffffffffff6f669dfd61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd1d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb211c",
    x"020900000000000002aa00000000000000fb336ad21c",
    x"030b00000000000002aafffffffffffff50003e8e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5fb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b8b1c",
    x"070a00000000000002aafffffffffffff8ef35f4521c",
    x"080200000000000002aafffffffffffff6f669dfd41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd191c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb221c",
    x"020900000000000002aa00000000000000fb336acc1c",
    x"030b00000000000002aafffffffffffff50003e8e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5f91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b851c",
    x"070a00000000000002aafffffffffffff8ef35f44f1c",
    x"080200000000000002aafffffffffffff6f669dfd11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd151c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb231c",
    x"020900000000000002aa00000000000000fb336ac71c",
    x"030b00000000000002aafffffffffffff50003e8ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5f61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b7f1c",
    x"070a00000000000002aafffffffffffff8ef35f44b1c",
    x"080200000000000002aafffffffffffff6f669dfcf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb241c",
    x"020900000000000002aa00000000000000fb336ac11c",
    x"030b00000000000002aafffffffffffff50003e8eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5f41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f381c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b791c",
    x"070a00000000000002aafffffffffffff8ef35f4471c",
    x"080200000000000002aafffffffffffff6f669dfcc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd0c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb251c",
    x"020900000000000002aa00000000000000fb336abb1c",
    x"030b00000000000002aafffffffffffff50003e8eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5f11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b731c",
    x"070a00000000000002aafffffffffffff8ef35f4441c",
    x"080200000000000002aafffffffffffff6f669dfca1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd081c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb261c",
    x"020900000000000002aa00000000000000fb336ab61c",
    x"030b00000000000002aafffffffffffff50003e8ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5ef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b6c1c",
    x"070a00000000000002aafffffffffffff8ef35f4401c",
    x"080200000000000002aafffffffffffff6f669dfc81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd041c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb271c",
    x"020900000000000002aa00000000000000fb336ab01c",
    x"030b00000000000002aafffffffffffff50003e8ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5ed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b661c",
    x"070a00000000000002aafffffffffffff8ef35f43c1c",
    x"080200000000000002aafffffffffffff6f669dfc51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cd001c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb291c",
    x"020900000000000002aa00000000000000fb336aaa1c",
    x"030b00000000000002aafffffffffffff50003e8ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5ea1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f380d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b601c",
    x"070a00000000000002aafffffffffffff8ef35f4391c",
    x"080200000000000002aafffffffffffff6f669dfc31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccfc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb2a1c",
    x"020900000000000002aa00000000000000fb336aa51c",
    x"030b00000000000002aafffffffffffff50003e8ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5e81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f380a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b5a1c",
    x"070a00000000000002aafffffffffffff8ef35f4351c",
    x"080200000000000002aafffffffffffff6f669dfc01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccf81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb2b1c",
    x"020900000000000002aa00000000000000fb336a9f1c",
    x"030b00000000000002aafffffffffffff50003e8f01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5e51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b541c",
    x"070a00000000000002aafffffffffffff8ef35f4311c",
    x"080200000000000002aafffffffffffff6f669dfbe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccf31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb2c1c",
    x"020900000000000002aa00000000000000fb336a9a1c",
    x"030b00000000000002aafffffffffffff50003e8f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5e31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f38031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b4e1c",
    x"070a00000000000002aafffffffffffff8ef35f42e1c",
    x"080200000000000002aafffffffffffff6f669dfbc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccef1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb2d1c",
    x"020900000000000002aa00000000000000fb336a941c",
    x"030b00000000000002aafffffffffffff50003e8f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5e01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b471c",
    x"070a00000000000002aafffffffffffff8ef35f42a1c",
    x"080200000000000002aafffffffffffff6f669dfb91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cceb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb2e1c",
    x"020900000000000002aa00000000000000fb336a8e1c",
    x"030b00000000000002aafffffffffffff50003e8f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5de1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b411c",
    x"070a00000000000002aafffffffffffff8ef35f4261c",
    x"080200000000000002aafffffffffffff6f669dfb71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266cce71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbeb2f1c",
    x"0209000000000000029a00000000000000fb336a891c",
    x"030b000000000000029afffffffffffff50003e8f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc5db1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f37f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd1b3b1c",
    x"070a000000000000029afffffffffffff8ef35f4221c",
    x"0802000000000000029afffffffffffff6f669dfb41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cce31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb301c",
    x"020900000000000002aa00000000000000fb336a831c",
    x"030b00000000000002aafffffffffffff50003e8f51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5d91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b351c",
    x"070a00000000000002aafffffffffffff8ef35f41f1c",
    x"080200000000000002aafffffffffffff6f669dfb21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266ccdf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb321c",
    x"0209000000000000031f00000000000000fb336a7e1c",
    x"030b000000000000031ffffffffffffff50003e8f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc5d61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f37f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1b2f1c",
    x"070a000000000000031ffffffffffffff8ef35f41b1c",
    x"0802000000000000031ffffffffffffff6f669dfaf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266ccda1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb331c",
    x"020900000000000000ae00000000000000fb336a781c",
    x"030b00000000000000aefffffffffffff50003e8f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc5d41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f37ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1b291c",
    x"070a00000000000000aefffffffffffff8ef35f4171c",
    x"080200000000000000aefffffffffffff6f669dfad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ccd61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb341c",
    x"020900000000000001a400000000000000fb336a721c",
    x"030b00000000000001a4fffffffffffff50003e8f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc5d11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f37e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1b221c",
    x"070a00000000000001a4fffffffffffff8ef35f4141c",
    x"080200000000000001a4fffffffffffff6f669dfab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266ccd21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbeb351c",
    x"0209000000000000029600000000000000fb336a6d1c",
    x"030b0000000000000296fffffffffffff50003e8f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dc5cf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f37e51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd1b1c1c",
    x"070a0000000000000296fffffffffffff8ef35f4101c",
    x"08020000000000000296fffffffffffff6f669dfa81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb361c",
    x"020900000000000002aa00000000000000fb336a671c",
    x"030b00000000000002aafffffffffffff50003e8f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b161c",
    x"070a00000000000002aafffffffffffff8ef35f40c1c",
    x"080200000000000002aafffffffffffff6f669dfa61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266ccca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbeb371c",
    x"020900000000000002a600000000000000fb336a621c",
    x"030b00000000000002a6fffffffffffff50003e8fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc5ca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f37de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd1b101c",
    x"070a00000000000002a6fffffffffffff8ef35f4091c",
    x"080200000000000002a6fffffffffffff6f669dfa31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccc61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb381c",
    x"020900000000000002aa00000000000000fb336a5c1c",
    x"030b00000000000002aafffffffffffff50003e8fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37db1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b0a1c",
    x"070a00000000000002aafffffffffffff8ef35f4051c",
    x"080200000000000002aafffffffffffff6f669dfa11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccc11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb391c",
    x"020900000000000002aa00000000000000fb336a561c",
    x"030b00000000000002aafffffffffffff50003e8fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37d71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1b041c",
    x"070a00000000000002aafffffffffffff8ef35f4011c",
    x"080200000000000002aafffffffffffff6f669df9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccbd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb3b1c",
    x"020900000000000002aa00000000000000fb336a511c",
    x"030b00000000000002aafffffffffffff50003e8fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37d31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1afd1c",
    x"070a00000000000002aafffffffffffff8ef35f3fe1c",
    x"080200000000000002aafffffffffffff6f669df9c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccb91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb3c1c",
    x"020900000000000002aa00000000000000fb336a4b1c",
    x"030b00000000000002aafffffffffffff50003e8fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5c01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37d01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1af71c",
    x"070a00000000000002aafffffffffffff8ef35f3fa1c",
    x"080200000000000002aafffffffffffff6f669df9a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccb51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb3d1c",
    x"020900000000000002aa00000000000000fb336a451c",
    x"030b00000000000002aafffffffffffff50003e8ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37cc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1af11c",
    x"070a00000000000002aafffffffffffff8ef35f3f61c",
    x"080200000000000002aafffffffffffff6f669df971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccb11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb3e1c",
    x"020900000000000002aa00000000000000fb336a401c",
    x"030b00000000000002aafffffffffffff50003e9001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37c81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1aeb1c",
    x"070a00000000000002aafffffffffffff8ef35f3f31c",
    x"080200000000000002aafffffffffffff6f669df951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ccad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb3f1c",
    x"020900000000000002aa00000000000000fb336a3a1c",
    x"030b00000000000002aafffffffffffff50003e9011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37c51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1ae51c",
    x"070a00000000000002aafffffffffffff8ef35f3ef1c",
    x"080200000000000002aafffffffffffff6f669df931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cca81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb401c",
    x"020900000000000002aa00000000000000fb336a351c",
    x"030b00000000000002aafffffffffffff50003e9021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37c11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1adf1c",
    x"070a00000000000002aafffffffffffff8ef35f3eb1c",
    x"080200000000000002aafffffffffffff6f669df901c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cca41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb411c",
    x"020900000000000002aa00000000000000fb336a2f1c",
    x"030b00000000000002aafffffffffffff50003e9031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1ad81c",
    x"070a00000000000002aafffffffffffff8ef35f3e71c",
    x"080200000000000002aafffffffffffff6f669df8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cca01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb421c",
    x"020900000000000002aa00000000000000fb336a291c",
    x"030b00000000000002aafffffffffffff50003e9031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5b11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37ba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1ad21c",
    x"070a00000000000002aafffffffffffff8ef35f3e41c",
    x"080200000000000002aafffffffffffff6f669df8b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cc9c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb441c",
    x"020900000000000002aa00000000000000fb336a241c",
    x"030b00000000000002aafffffffffffff50003e9041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37b61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1acc1c",
    x"070a00000000000002aafffffffffffff8ef35f3e01c",
    x"080200000000000002aafffffffffffff6f669df891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cc981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb451c",
    x"020900000000000002aa00000000000000fb336a1e1c",
    x"030b00000000000002aafffffffffffff50003e9051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5ac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1ac61c",
    x"070a00000000000002aafffffffffffff8ef35f3dc1c",
    x"080200000000000002aafffffffffffff6f669df871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266cc941c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbeb461c",
    x"0209000000000000029a00000000000000fb336a191c",
    x"030b000000000000029afffffffffffff50003e9061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc5aa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f37af1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd1ac01c",
    x"070a000000000000029afffffffffffff8ef35f3d91c",
    x"0802000000000000029afffffffffffff6f669df841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cc8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb471c",
    x"020900000000000002aa00000000000000fb336a131c",
    x"030b00000000000002aafffffffffffff50003e9071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5a71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37ab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1ab91c",
    x"070a00000000000002aafffffffffffff8ef35f3d51c",
    x"080200000000000002aafffffffffffff6f669df821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cc8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb481c",
    x"0209000000000000031f00000000000000fb336a0d1c",
    x"030b000000000000031ffffffffffffff50003e9081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc5a51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f37a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1ab31c",
    x"070a000000000000031ffffffffffffff8ef35f3d11c",
    x"0802000000000000031ffffffffffffff6f669df7f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cc871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb491c",
    x"020900000000000000ae00000000000000fb336a081c",
    x"030b00000000000000aefffffffffffff50003e9091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc5a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f37a41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1aad1c",
    x"070a00000000000000aefffffffffffff8ef35f3ce1c",
    x"080200000000000000aefffffffffffff6f669df7d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cc831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb4a1c",
    x"020900000000000001a400000000000000fb336a021c",
    x"030b00000000000001a4fffffffffffff50003e90a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc5a01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f37a01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1aa71c",
    x"070a00000000000001a4fffffffffffff8ef35f3ca1c",
    x"080200000000000001a4fffffffffffff6f669df7a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266cc7f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbeb4b1c",
    x"0209000000000000019600000000000000fb3369fd1c",
    x"030b0000000000000196fffffffffffff50003e90b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc59d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f379d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001960000000000000004cd1aa11c",
    x"070a0000000000000196fffffffffffff8ef35f3c61c",
    x"08020000000000000196fffffffffffff6f669df781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc7b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb4d1c",
    x"0209000000000000015500000000000000fb3369f71c",
    x"030b0000000000000155fffffffffffff50003e90c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc59b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37991c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a9b1c",
    x"070a0000000000000155fffffffffffff8ef35f3c31c",
    x"08020000000000000155fffffffffffff6f669df761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb4e1c",
    x"0209000000000000015500000000000000fb3369f11c",
    x"030b0000000000000155fffffffffffff50003e90d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a941c",
    x"070a0000000000000155fffffffffffff8ef35f3bf1c",
    x"08020000000000000155fffffffffffff6f669df731c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb4f1c",
    x"0209000000000000015500000000000000fb3369ec1c",
    x"030b0000000000000155fffffffffffff50003e90e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a8e1c",
    x"070a0000000000000155fffffffffffff8ef35f3bb1c",
    x"08020000000000000155fffffffffffff6f669df711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc6e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb501c",
    x"0209000000000000015500000000000000fb3369e61c",
    x"030b0000000000000155fffffffffffff50003e90e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f378e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a881c",
    x"070a0000000000000155fffffffffffff8ef35f3b81c",
    x"08020000000000000155fffffffffffff6f669df6e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc6a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb511c",
    x"0209000000000000015500000000000000fb3369e01c",
    x"030b0000000000000155fffffffffffff50003e90f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f378b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a821c",
    x"070a0000000000000155fffffffffffff8ef35f3b41c",
    x"08020000000000000155fffffffffffff6f669df6c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb521c",
    x"0209000000000000015500000000000000fb3369db1c",
    x"030b0000000000000155fffffffffffff50003e9101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc58e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37871c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a7c1c",
    x"070a0000000000000155fffffffffffff8ef35f3b01c",
    x"08020000000000000155fffffffffffff6f669df6a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb531c",
    x"0209000000000000015500000000000000fb3369d51c",
    x"030b0000000000000155fffffffffffff50003e9111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc58c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37831c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a761c",
    x"070a0000000000000155fffffffffffff8ef35f3ac1c",
    x"08020000000000000155fffffffffffff6f669df671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb541c",
    x"0209000000000000015500000000000000fb3369d01c",
    x"030b0000000000000155fffffffffffff50003e9121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a6f1c",
    x"070a0000000000000155fffffffffffff8ef35f3a91c",
    x"08020000000000000155fffffffffffff6f669df651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb561c",
    x"0209000000000000015500000000000000fb3369ca1c",
    x"030b0000000000000155fffffffffffff50003e9131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f377c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a691c",
    x"070a0000000000000155fffffffffffff8ef35f3a51c",
    x"08020000000000000155fffffffffffff6f669df621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb571c",
    x"0209000000000000015500000000000000fb3369c41c",
    x"030b0000000000000155fffffffffffff50003e9141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a631c",
    x"070a0000000000000155fffffffffffff8ef35f3a11c",
    x"08020000000000000155fffffffffffff6f669df601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb581c",
    x"0209000000000000015500000000000000fb3369bf1c",
    x"030b0000000000000155fffffffffffff50003e9151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37751c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a5d1c",
    x"070a0000000000000155fffffffffffff8ef35f39e1c",
    x"08020000000000000155fffffffffffff6f669df5e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc4d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb591c",
    x"0209000000000000015500000000000000fb3369b91c",
    x"030b0000000000000155fffffffffffff50003e9161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc57f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a571c",
    x"070a0000000000000155fffffffffffff8ef35f39a1c",
    x"08020000000000000155fffffffffffff6f669df5b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb5a1c",
    x"0209000000000000015500000000000000fb3369b41c",
    x"030b0000000000000155fffffffffffff50003e9171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc57d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f376e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a511c",
    x"070a0000000000000155fffffffffffff8ef35f3961c",
    x"08020000000000000155fffffffffffff6f669df591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb5b1c",
    x"0209000000000000015500000000000000fb3369ae1c",
    x"030b0000000000000155fffffffffffff50003e9181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc57a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f376a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a4a1c",
    x"070a0000000000000155fffffffffffff8ef35f3931c",
    x"08020000000000000155fffffffffffff6f669df561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266cc401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbeb5c1c",
    x"020900000000000002a500000000000000fb3369a81c",
    x"030b00000000000002a5fffffffffffff50003e9191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc5781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f37661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd1a441c",
    x"070a00000000000002a5fffffffffffff8ef35f38f1c",
    x"080200000000000002a5fffffffffffff6f669df541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cc3c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb5e1c",
    x"020900000000000002aa00000000000000fb3369a31c",
    x"030b00000000000002aafffffffffffff50003e91a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37631c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1a3e1c",
    x"070a00000000000002aafffffffffffff8ef35f38b1c",
    x"080200000000000002aafffffffffffff6f669df521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cc381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb5f1c",
    x"0209000000000000031f00000000000000fb33699d1c",
    x"030b000000000000031ffffffffffffff50003e91a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc5731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f375f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd1a381c",
    x"070a000000000000031ffffffffffffff8ef35f3881c",
    x"0802000000000000031ffffffffffffff6f669df4f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cc341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb601c",
    x"020900000000000000ae00000000000000fb3369971c",
    x"030b00000000000000aefffffffffffff50003e91b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc5701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f375c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd1a321c",
    x"070a00000000000000aefffffffffffff8ef35f3841c",
    x"080200000000000000aefffffffffffff6f669df4d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cc2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb611c",
    x"020900000000000001a400000000000000fb3369921c",
    x"030b00000000000001a4fffffffffffff50003e91c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc56e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f37581c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd1a2b1c",
    x"070a00000000000001a4fffffffffffff8ef35f3801c",
    x"080200000000000001a4fffffffffffff6f669df4a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266cc2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbeb621c",
    x"020900000000000002a600000000000000fb33698c1c",
    x"030b00000000000002a6fffffffffffff50003e91d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc56b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f37541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd1a251c",
    x"070a00000000000002a6fffffffffffff8ef35f37c1c",
    x"080200000000000002a6fffffffffffff6f669df481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cc271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb631c",
    x"020900000000000002aa00000000000000fb3369871c",
    x"030b00000000000002aafffffffffffff50003e91e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f37511c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd1a1f1c",
    x"070a00000000000002aafffffffffffff8ef35f3791c",
    x"080200000000000002aafffffffffffff6f669df451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266cc231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbeb641c",
    x"0209000000000000015600000000000000fb3369811c",
    x"030b0000000000000156fffffffffffff50003e91f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc5661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f374d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd1a191c",
    x"070a0000000000000156fffffffffffff8ef35f3751c",
    x"08020000000000000156fffffffffffff6f669df431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc1f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb651c",
    x"0209000000000000015500000000000000fb33697b1c",
    x"030b0000000000000155fffffffffffff50003e9201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a131c",
    x"070a0000000000000155fffffffffffff8ef35f3711c",
    x"08020000000000000155fffffffffffff6f669df411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc1b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb671c",
    x"0209000000000000015500000000000000fb3369761c",
    x"030b0000000000000155fffffffffffff50003e9211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37461c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a0d1c",
    x"070a0000000000000155fffffffffffff8ef35f36e1c",
    x"08020000000000000155fffffffffffff6f669df3e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb681c",
    x"0209000000000000015500000000000000fb3369701c",
    x"030b0000000000000155fffffffffffff50003e9221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc55f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a061c",
    x"070a0000000000000155fffffffffffff8ef35f36a1c",
    x"08020000000000000155fffffffffffff6f669df3c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb691c",
    x"0209000000000000015500000000000000fb33696b1c",
    x"030b0000000000000155fffffffffffff50003e9231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc55c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f373f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd1a001c",
    x"070a0000000000000155fffffffffffff8ef35f3661c",
    x"08020000000000000155fffffffffffff6f669df391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc0e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb6a1c",
    x"0209000000000000015500000000000000fb3369651c",
    x"030b0000000000000155fffffffffffff50003e9241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc55a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f373b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19fa1c",
    x"070a0000000000000155fffffffffffff8ef35f3631c",
    x"08020000000000000155fffffffffffff6f669df371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc0a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb6b1c",
    x"0209000000000000015500000000000000fb33695f1c",
    x"030b0000000000000155fffffffffffff50003e9251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19f41c",
    x"070a0000000000000155fffffffffffff8ef35f35f1c",
    x"08020000000000000155fffffffffffff6f669df351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb6c1c",
    x"0209000000000000015500000000000000fb33695a1c",
    x"030b0000000000000155fffffffffffff50003e9251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19ee1c",
    x"070a0000000000000155fffffffffffff8ef35f35b1c",
    x"08020000000000000155fffffffffffff6f669df321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cc021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb6d1c",
    x"0209000000000000015500000000000000fb3369541c",
    x"030b0000000000000155fffffffffffff50003e9261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37301c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19e81c",
    x"070a0000000000000155fffffffffffff8ef35f3581c",
    x"08020000000000000155fffffffffffff6f669df301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbfd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb6e1c",
    x"0209000000000000015500000000000000fb33694f1c",
    x"030b0000000000000155fffffffffffff50003e9271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f372c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19e11c",
    x"070a0000000000000155fffffffffffff8ef35f3541c",
    x"08020000000000000155fffffffffffff6f669df2d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbf91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb701c",
    x"0209000000000000015500000000000000fb3369491c",
    x"030b0000000000000155fffffffffffff50003e9281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc54e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19db1c",
    x"070a0000000000000155fffffffffffff8ef35f3501c",
    x"08020000000000000155fffffffffffff6f669df2b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbf51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb711c",
    x"0209000000000000015500000000000000fb3369431c",
    x"030b0000000000000155fffffffffffff50003e9291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc54b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37251c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19d51c",
    x"070a0000000000000155fffffffffffff8ef35f34c1c",
    x"08020000000000000155fffffffffffff6f669df291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbf11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb721c",
    x"0209000000000000015500000000000000fb33693e1c",
    x"030b0000000000000155fffffffffffff50003e92a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37221c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19cf1c",
    x"070a0000000000000155fffffffffffff8ef35f3491c",
    x"08020000000000000155fffffffffffff6f669df261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266cbed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbeb731c",
    x"0209000000000000016500000000000000fb3369381c",
    x"030b0000000000000165fffffffffffff50003e92b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc5461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f371e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd19c91c",
    x"070a0000000000000165fffffffffffff8ef35f3451c",
    x"08020000000000000165fffffffffffff6f669df241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cbe91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb741c",
    x"020900000000000002aa00000000000000fb3369321c",
    x"030b00000000000002aafffffffffffff50003e92c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f371a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd19c31c",
    x"070a00000000000002aafffffffffffff8ef35f3411c",
    x"080200000000000002aafffffffffffff6f669df211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cbe41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb751c",
    x"0209000000000000031f00000000000000fb33692d1c",
    x"030b000000000000031ffffffffffffff50003e92d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc5411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f37171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd19bc1c",
    x"070a000000000000031ffffffffffffff8ef35f33e1c",
    x"0802000000000000031ffffffffffffff6f669df1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cbe01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb761c",
    x"020900000000000000ae00000000000000fb3369271c",
    x"030b00000000000000aefffffffffffff50003e92e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc53f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f37131c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd19b61c",
    x"070a00000000000000aefffffffffffff8ef35f33a1c",
    x"080200000000000000aefffffffffffff6f669df1d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cbdc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb771c",
    x"020900000000000001a400000000000000fb3369221c",
    x"030b00000000000001a4fffffffffffff50003e92f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc53c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f370f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd19b01c",
    x"070a00000000000001a4fffffffffffff8ef35f3361c",
    x"080200000000000001a4fffffffffffff6f669df1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266cbd81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbeb791c",
    x"020900000000000001a600000000000000fb33691c1c",
    x"030b00000000000001a6fffffffffffff50003e9301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc53a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f370c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd19aa1c",
    x"070a00000000000001a6fffffffffffff8ef35f3331c",
    x"080200000000000001a6fffffffffffff6f669df181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbd41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb7a1c",
    x"0209000000000000015500000000000000fb3369161c",
    x"030b0000000000000155fffffffffffff50003e9301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37081c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19a41c",
    x"070a0000000000000155fffffffffffff8ef35f32f1c",
    x"08020000000000000155fffffffffffff6f669df151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbd01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb7b1c",
    x"0209000000000000015500000000000000fb3369111c",
    x"030b0000000000000155fffffffffffff50003e9311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5351c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd199d1c",
    x"070a0000000000000155fffffffffffff8ef35f32b1c",
    x"08020000000000000155fffffffffffff6f669df131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbcb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb7c1c",
    x"0209000000000000015500000000000000fb33690b1c",
    x"030b0000000000000155fffffffffffff50003e9321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f37011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19971c",
    x"070a0000000000000155fffffffffffff8ef35f3281c",
    x"08020000000000000155fffffffffffff6f669df101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbc71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb7d1c",
    x"0209000000000000015500000000000000fb3369061c",
    x"030b0000000000000155fffffffffffff50003e9331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5301c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36fd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19911c",
    x"070a0000000000000155fffffffffffff8ef35f3241c",
    x"08020000000000000155fffffffffffff6f669df0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbc31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb7e1c",
    x"0209000000000000015500000000000000fb3369001c",
    x"030b0000000000000155fffffffffffff50003e9341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc52d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36fa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd198b1c",
    x"070a0000000000000155fffffffffffff8ef35f3201c",
    x"08020000000000000155fffffffffffff6f669df0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbbf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb7f1c",
    x"0209000000000000015500000000000000fb3368fa1c",
    x"030b0000000000000155fffffffffffff50003e9351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc52b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36f61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19851c",
    x"070a0000000000000155fffffffffffff8ef35f31c1c",
    x"08020000000000000155fffffffffffff6f669df091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbbb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb811c",
    x"0209000000000000015500000000000000fb3368f51c",
    x"030b0000000000000155fffffffffffff50003e9361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36f21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd197f1c",
    x"070a0000000000000155fffffffffffff8ef35f3191c",
    x"08020000000000000155fffffffffffff6f669df071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbb71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb821c",
    x"0209000000000000015500000000000000fb3368ef1c",
    x"030b0000000000000155fffffffffffff50003e9371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36ef1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19781c",
    x"070a0000000000000155fffffffffffff8ef35f3151c",
    x"08020000000000000155fffffffffffff6f669df041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbb21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb831c",
    x"0209000000000000015500000000000000fb3368e91c",
    x"030b0000000000000155fffffffffffff50003e9381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36eb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19721c",
    x"070a0000000000000155fffffffffffff8ef35f3111c",
    x"08020000000000000155fffffffffffff6f669df021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb841c",
    x"0209000000000000015500000000000000fb3368e41c",
    x"030b0000000000000155fffffffffffff50003e9391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36e81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd196c1c",
    x"070a0000000000000155fffffffffffff8ef35f30e1c",
    x"08020000000000000155fffffffffffff6f669df001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cbaa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb851c",
    x"0209000000000000015500000000000000fb3368de1c",
    x"030b0000000000000155fffffffffffff50003e93a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc51e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36e41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19661c",
    x"070a0000000000000155fffffffffffff8ef35f30a1c",
    x"08020000000000000155fffffffffffff6f669defd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cba61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb861c",
    x"0209000000000000015500000000000000fb3368d91c",
    x"030b0000000000000155fffffffffffff50003e93b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc51c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36e01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19601c",
    x"070a0000000000000155fffffffffffff8ef35f3061c",
    x"08020000000000000155fffffffffffff6f669defb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cba21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb871c",
    x"0209000000000000015500000000000000fb3368d31c",
    x"030b0000000000000155fffffffffffff50003e93b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36dd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd195a1c",
    x"070a0000000000000155fffffffffffff8ef35f3031c",
    x"08020000000000000155fffffffffffff6f669def81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb9e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb881c",
    x"0209000000000000015500000000000000fb3368cd1c",
    x"030b0000000000000155fffffffffffff50003e93c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19531c",
    x"070a0000000000000155fffffffffffff8ef35f2ff1c",
    x"08020000000000000155fffffffffffff6f669def61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cb991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbeb8a1c",
    x"0209000000000000029500000000000000fb3368c81c",
    x"030b0000000000000295fffffffffffff50003e93d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc5141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f36d51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd194d1c",
    x"070a0000000000000295fffffffffffff8ef35f2fb1c",
    x"08020000000000000295fffffffffffff6f669def41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeb8b1c",
    x"020900000000000002aa00000000000000fb3368c21c",
    x"030b00000000000002aafffffffffffff50003e93e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc5121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36d21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd19471c",
    x"070a00000000000002aafffffffffffff8ef35f2f81c",
    x"080200000000000002aafffffffffffff6f669def11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cb911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeb8c1c",
    x"0209000000000000031f00000000000000fb3368bd1c",
    x"030b000000000000031ffffffffffffff50003e93f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc50f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f36ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd19411c",
    x"070a000000000000031ffffffffffffff8ef35f2f41c",
    x"0802000000000000031ffffffffffffff6f669deef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cb8d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeb8d1c",
    x"020900000000000000ae00000000000000fb3368b71c",
    x"030b00000000000000aefffffffffffff50003e9401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc50d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f36cb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd193b1c",
    x"070a00000000000000aefffffffffffff8ef35f2f01c",
    x"080200000000000000aefffffffffffff6f669deec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cb891c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeb8e1c",
    x"020900000000000001a400000000000000fb3368b11c",
    x"030b00000000000001a4fffffffffffff50003e9411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc50a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f36c71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd19341c",
    x"070a00000000000001a4fffffffffffff8ef35f2ec1c",
    x"080200000000000001a4fffffffffffff6f669deea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266cb851c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbeb8f1c",
    x"0209000000000000016600000000000000fb3368ac1c",
    x"030b0000000000000166fffffffffffff50003e9421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc5081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f36c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd192e1c",
    x"070a0000000000000166fffffffffffff8ef35f2e91c",
    x"08020000000000000166fffffffffffff6f669dee71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb901c",
    x"0209000000000000015500000000000000fb3368a61c",
    x"030b0000000000000155fffffffffffff50003e9431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36c01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19281c",
    x"070a0000000000000155fffffffffffff8ef35f2e51c",
    x"08020000000000000155fffffffffffff6f669dee51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb7c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb911c",
    x"0209000000000000015500000000000000fb3368a11c",
    x"030b0000000000000155fffffffffffff50003e9441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36bc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19221c",
    x"070a0000000000000155fffffffffffff8ef35f2e11c",
    x"08020000000000000155fffffffffffff6f669dee31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb931c",
    x"0209000000000000015500000000000000fb33689b1c",
    x"030b0000000000000155fffffffffffff50003e9451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc5001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36b81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd191c1c",
    x"070a0000000000000155fffffffffffff8ef35f2de1c",
    x"08020000000000000155fffffffffffff6f669dee01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb741c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb941c",
    x"0209000000000000015500000000000000fb3368951c",
    x"030b0000000000000155fffffffffffff50003e9461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4fe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36b51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19161c",
    x"070a0000000000000155fffffffffffff8ef35f2da1c",
    x"08020000000000000155fffffffffffff6f669dede1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb701c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb951c",
    x"0209000000000000015500000000000000fb3368901c",
    x"030b0000000000000155fffffffffffff50003e9461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4fb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36b11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd190f1c",
    x"070a0000000000000155fffffffffffff8ef35f2d61c",
    x"08020000000000000155fffffffffffff6f669dedb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb6c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb961c",
    x"0209000000000000015500000000000000fb33688a1c",
    x"030b0000000000000155fffffffffffff50003e9471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4f91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36ae1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19091c",
    x"070a0000000000000155fffffffffffff8ef35f2d31c",
    x"08020000000000000155fffffffffffff6f669ded91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb971c",
    x"0209000000000000015500000000000000fb3368841c",
    x"030b0000000000000155fffffffffffff50003e9481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4f61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36aa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd19031c",
    x"070a0000000000000155fffffffffffff8ef35f2cf1c",
    x"08020000000000000155fffffffffffff6f669ded71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb981c",
    x"0209000000000000015500000000000000fb33687f1c",
    x"030b0000000000000155fffffffffffff50003e9491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4f41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36a61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18fd1c",
    x"070a0000000000000155fffffffffffff8ef35f2cb1c",
    x"08020000000000000155fffffffffffff6f669ded41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb5f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb991c",
    x"0209000000000000015500000000000000fb3368791c",
    x"030b0000000000000155fffffffffffff50003e94a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4f11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36a31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18f71c",
    x"070a0000000000000155fffffffffffff8ef35f2c71c",
    x"08020000000000000155fffffffffffff6f669ded21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb5b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb9a1c",
    x"0209000000000000015500000000000000fb3368741c",
    x"030b0000000000000155fffffffffffff50003e94b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4ef1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f369f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18f11c",
    x"070a0000000000000155fffffffffffff8ef35f2c41c",
    x"08020000000000000155fffffffffffff6f669decf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb571c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb9c1c",
    x"0209000000000000015500000000000000fb33686e1c",
    x"030b0000000000000155fffffffffffff50003e94c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4ec1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f369b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18ea1c",
    x"070a0000000000000155fffffffffffff8ef35f2c01c",
    x"08020000000000000155fffffffffffff6f669decd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb531c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb9d1c",
    x"0209000000000000015500000000000000fb3368681c",
    x"030b0000000000000155fffffffffffff50003e94d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4ea1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18e41c",
    x"070a0000000000000155fffffffffffff8ef35f2bc1c",
    x"08020000000000000155fffffffffffff6f669decb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb4e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb9e1c",
    x"0209000000000000015500000000000000fb3368631c",
    x"030b0000000000000155fffffffffffff50003e94e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4e71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18de1c",
    x"070a0000000000000155fffffffffffff8ef35f2b91c",
    x"08020000000000000155fffffffffffff6f669dec81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb4a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeb9f1c",
    x"0209000000000000015500000000000000fb33685d1c",
    x"030b0000000000000155fffffffffffff50003e94f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4e51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18d81c",
    x"070a0000000000000155fffffffffffff8ef35f2b51c",
    x"08020000000000000155fffffffffffff6f669dec61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266cb461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbeba01c",
    x"0209000000000000016500000000000000fb3368581c",
    x"030b0000000000000165fffffffffffff50003e9501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc4e21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f368d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd18d21c",
    x"070a0000000000000165fffffffffffff8ef35f2b11c",
    x"08020000000000000165fffffffffffff6f669dec31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266cb421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeba11c",
    x"0209000000000000015500000000000000fb3368521c",
    x"030b0000000000000155fffffffffffff50003e9501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4e01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd18cc1c",
    x"070a0000000000000155fffffffffffff8ef35f2ae1c",
    x"08020000000000000155fffffffffffff6f669dec11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266cb3e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeba21c",
    x"0209000000000000031f00000000000000fb33684c1c",
    x"030b000000000000031ffffffffffffff50003e9511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc4de1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f36861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd18c51c",
    x"070a000000000000031ffffffffffffff8ef35f2aa1c",
    x"0802000000000000031ffffffffffffff6f669debe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cb3a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeba41c",
    x"020900000000000000ae00000000000000fb3368471c",
    x"030b00000000000000aefffffffffffff50003e9521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc4db1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f36821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd18bf1c",
    x"070a00000000000000aefffffffffffff8ef35f2a61c",
    x"080200000000000000aefffffffffffff6f669debc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cb351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeba51c",
    x"020900000000000001a400000000000000fb3368411c",
    x"030b00000000000001a4fffffffffffff50003e9531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc4d91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f367e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd18b91c",
    x"070a00000000000001a4fffffffffffff8ef35f2a31c",
    x"080200000000000001a4fffffffffffff6f669deba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266cb311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbeba61c",
    x"0209000000000000026600000000000000fb33683b1c",
    x"030b0000000000000266fffffffffffff50003e9541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc4d61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f367b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002660000000000000004cd18b31c",
    x"070a0000000000000266fffffffffffff8ef35f29f1c",
    x"08020000000000000266fffffffffffff6f669deb71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb2d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeba71c",
    x"020900000000000002aa00000000000000fb3368361c",
    x"030b00000000000002aafffffffffffff50003e9551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4d41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18ad1c",
    x"070a00000000000002aafffffffffffff8ef35f29b1c",
    x"080200000000000002aafffffffffffff6f669deb51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb291c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeba81c",
    x"020900000000000002aa00000000000000fb3368301c",
    x"030b00000000000002aafffffffffffff50003e9561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4d11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18a61c",
    x"070a00000000000002aafffffffffffff8ef35f2971c",
    x"080200000000000002aafffffffffffff6f669deb21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb251c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbeba91c",
    x"020900000000000002aa00000000000000fb33682b1c",
    x"030b00000000000002aafffffffffffff50003e9571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4cf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36701c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18a01c",
    x"070a00000000000002aafffffffffffff8ef35f2941c",
    x"080200000000000002aafffffffffffff6f669deb01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebaa1c",
    x"020900000000000002aa00000000000000fb3368251c",
    x"030b00000000000002aafffffffffffff50003e9581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f366c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd189a1c",
    x"070a00000000000002aafffffffffffff8ef35f2901c",
    x"080200000000000002aafffffffffffff6f669deae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb1c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebab1c",
    x"020900000000000002aa00000000000000fb33681f1c",
    x"030b00000000000002aafffffffffffff50003e9591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4ca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18941c",
    x"070a00000000000002aafffffffffffff8ef35f28c1c",
    x"080200000000000002aafffffffffffff6f669deab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebad1c",
    x"020900000000000002aa00000000000000fb33681a1c",
    x"030b00000000000002aafffffffffffff50003e95a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd188e1c",
    x"070a00000000000002aafffffffffffff8ef35f2891c",
    x"080200000000000002aafffffffffffff6f669dea91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebae1c",
    x"020900000000000002aa00000000000000fb3368141c",
    x"030b00000000000002aafffffffffffff50003e95b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18881c",
    x"070a00000000000002aafffffffffffff8ef35f2851c",
    x"080200000000000002aafffffffffffff6f669dea61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebaf1c",
    x"020900000000000002aa00000000000000fb33680f1c",
    x"030b00000000000002aafffffffffffff50003e95b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f365e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18811c",
    x"070a00000000000002aafffffffffffff8ef35f2811c",
    x"080200000000000002aafffffffffffff6f669dea41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb0c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb01c",
    x"020900000000000002aa00000000000000fb3368091c",
    x"030b00000000000002aafffffffffffff50003e95c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4c01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f365a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd187b1c",
    x"070a00000000000002aafffffffffffff8ef35f27e1c",
    x"080200000000000002aafffffffffffff6f669dea21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb081c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb11c",
    x"020900000000000002aa00000000000000fb3368031c",
    x"030b00000000000002aafffffffffffff50003e95d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18751c",
    x"070a00000000000002aafffffffffffff8ef35f27a1c",
    x"080200000000000002aafffffffffffff6f669de9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cb031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb21c",
    x"020900000000000002aa00000000000000fb3367fe1c",
    x"030b00000000000002aafffffffffffff50003e95e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd186f1c",
    x"070a00000000000002aafffffffffffff8ef35f2761c",
    x"080200000000000002aafffffffffffff6f669de9d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266caff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb31c",
    x"020900000000000002aa00000000000000fb3367f81c",
    x"030b00000000000002aafffffffffffff50003e95f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f364f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18691c",
    x"070a00000000000002aafffffffffffff8ef35f2721c",
    x"080200000000000002aafffffffffffff6f669de9a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266cafb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb41c",
    x"020900000000000002aa00000000000000fb3367f21c",
    x"030b00000000000002aafffffffffffff50003e9601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f364c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18631c",
    x"070a00000000000002aafffffffffffff8ef35f26f1c",
    x"080200000000000002aafffffffffffff6f669de981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266caf71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb61c",
    x"020900000000000002aa00000000000000fb3367ed1c",
    x"030b00000000000002aafffffffffffff50003e9611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd185c1c",
    x"070a00000000000002aafffffffffffff8ef35f26b1c",
    x"080200000000000002aafffffffffffff6f669de961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266caf31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb71c",
    x"020900000000000002aa00000000000000fb3367e71c",
    x"030b00000000000002aafffffffffffff50003e9621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4b11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18561c",
    x"070a00000000000002aafffffffffffff8ef35f2671c",
    x"080200000000000002aafffffffffffff6f669de931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266caef1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebb81c",
    x"020900000000000002aa00000000000000fb3367e21c",
    x"030b00000000000002aafffffffffffff50003e9631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f36411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd18501c",
    x"070a00000000000002aafffffffffffff8ef35f2641c",
    x"080200000000000002aafffffffffffff6f669de911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266caea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbebb91c",
    x"0209000000000000031f00000000000000fb3367dc1c",
    x"030b000000000000031ffffffffffffff50003e9641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc4ac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f363d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd184a1c",
    x"070a000000000000031ffffffffffffff8ef35f2601c",
    x"0802000000000000031ffffffffffffff6f669de8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266cae61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbebba1c",
    x"020900000000000000ae00000000000000fb3367d61c",
    x"030b00000000000000aefffffffffffff50003e9651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc4a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f363a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd18441c",
    x"070a00000000000000aefffffffffffff8ef35f25c1c",
    x"080200000000000000aefffffffffffff6f669de8c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266cae21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbebbb1c",
    x"020900000000000001a400000000000000fb3367d11c",
    x"030b00000000000001a4fffffffffffff50003e9651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc4a71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f36361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd183d1c",
    x"070a00000000000001a4fffffffffffff8ef35f2591c",
    x"080200000000000001a4fffffffffffff6f669de891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266cade1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbebbc1c",
    x"020900000000000001aa00000000000000fb3367cb1c",
    x"030b00000000000001aafffffffffffff50003e9661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc4a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f36321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd18371c",
    x"070a00000000000001aafffffffffffff8ef35f2551c",
    x"080200000000000001aafffffffffffff6f669de871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cada1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbebbe1c",
    x"0209000000000000029500000000000000fb3367c61c",
    x"030b0000000000000295fffffffffffff50003e9671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc4a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f362f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd18311c",
    x"070a0000000000000295fffffffffffff8ef35f2511c",
    x"08020000000000000295fffffffffffff6f669de851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266cad61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbebbf1c",
    x"0209000000000000015a00000000000000fb3367c01c",
    x"030b000000000000015afffffffffffff50003e9681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc49f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f362b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd182b1c",
    x"070a000000000000015afffffffffffff8ef35f24d1c",
    x"0802000000000000015afffffffffffff6f669de821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266cad11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbebc01c",
    x"0209000000000000029500000000000000fb3367ba1c",
    x"030b0000000000000295fffffffffffff50003e9691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc49d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f36281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd18251c",
    x"070a0000000000000295fffffffffffff8ef35f24a1c",
    x"08020000000000000295fffffffffffff6f669de801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266cacd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbebc11c",
    x"020900000000000002a900000000000000fb3367b51c",
    x"030b0000000000000155fffffffffffff50003e96a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc49a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f36241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd181f1c",
    x"070a0000000000000155fffffffffffff8ef35f2461c",
    x"080200000000000002a9fffffffffffff6f669de7d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266cac91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebc21c",
    x"0209000000000000029a00000000000000fb3367af1c",
    x"030b0000000000000265fffffffffffff50003e96b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc4981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f36201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd18181c",
    x"070a0000000000000255fffffffffffff8ef35f2421c",
    x"080200000000000002a9fffffffffffff6f669de7b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266cac51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbebc31c",
    x"0209000000000000015a00000000000000fb3367aa1c",
    x"030b0000000000000265fffffffffffff50003e96c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc4951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f361d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd18121c",
    x"070a000000000000029afffffffffffff8ef35f23f1c",
    x"0802000000000000019afffffffffffff6f669de791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266cac11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbebc41c",
    x"0209000000000000019900000000000000fb3367a41c",
    x"030b0000000000000166fffffffffffff50003e96d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc4931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f36191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd180c1c",
    x"070a00000000000001a9fffffffffffff8ef35f23b1c",
    x"0802000000000000026afffffffffffff6f669de761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266cabd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002690000000000000b0bfbebc51c",
    x"0209000000000000016600000000000000fb33679e1c",
    x"030b00000000000001a6fffffffffffff50003e96e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc4901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f36151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd18061c",
    x"070a0000000000000199fffffffffffff8ef35f2371c",
    x"0802000000000000025afffffffffffff6f669de741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266cab81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebc71c",
    x"0209000000000000015500000000000000fb3367991c",
    x"030b000000000000015afffffffffffff50003e96f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc48e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f36121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd18001c",
    x"070a000000000000016afffffffffffff8ef35f2341c",
    x"0802000000000000025afffffffffffff6f669de711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266cab41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbebc81c",
    x"0209000000000000015a00000000000000fb3367931c",
    x"030b0000000000000295fffffffffffff50003e96f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc48b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f360e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd17fa1c",
    x"070a00000000000001aafffffffffffff8ef35f2301c",
    x"08020000000000000296fffffffffffff6f669de6f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266cab01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002990000000000000b0bfbebc91c",
    x"020900000000000001a900000000000000fb33678d1c",
    x"030b0000000000000299fffffffffffff50003e9701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dc4891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f360b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd17f31c",
    x"070a0000000000000165fffffffffffff8ef35f22c1c",
    x"0802000000000000016afffffffffffff6f669de6c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266caac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbebca1c",
    x"020900000000000002aa00000000000000fb3367881c",
    x"030b0000000000000169fffffffffffff50003e9711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc4861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f36071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd17ed1c",
    x"070a00000000000002a9fffffffffffff8ef35f2281c",
    x"08020000000000000199fffffffffffff6f669de6a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000299ffffffffffffff0266caa81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbebcb1c",
    x"0209000000000000029a00000000000000fb3367821c",
    x"030b000000000000019afffffffffffff50003e9721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc4841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f36031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd17e71c",
    x"070a000000000000016afffffffffffff8ef35f2251c",
    x"08020000000000000165fffffffffffff6f669de681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266caa41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbebcc1c",
    x"020900000000000002a600000000000000fb33677d1c",
    x"030b000000000000015afffffffffffff50003e9731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc4811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f36001c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd17e11c",
    x"070a000000000000025afffffffffffff8ef35f2211c",
    x"0802000000000000025afffffffffffff6f669de651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266ca9f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbebcd1c",
    x"0209000000000000029a00000000000000fb3367771c",
    x"030b0000000000000255fffffffffffff50003e9741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc47f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f35fc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd17db1c",
    x"070a0000000000000169fffffffffffff8ef35f21d1c",
    x"08020000000000000199fffffffffffff6f669de631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266ca9b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbebce1c",
    x"0209000000000000015900000000000000fb3367711c",
    x"030b00000000000002a6fffffffffffff50003e9751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc47c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd17d41c",
    x"070a00000000000002a6fffffffffffff8ef35f21a1c",
    x"0802000000000000016afffffffffffff6f669de601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266ca971c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbebd01c",
    x"0209000000000000031f00000000000000fb33676c1c",
    x"030b000000000000031ffffffffffffff50003e9761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc47a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f35f51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd17ce1c",
    x"070a000000000000031ffffffffffffff8ef35f2161c",
    x"0802000000000000031ffffffffffffff6f669de5e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266ca931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbebd11c",
    x"020900000000000000ae00000000000000fb3367661c",
    x"030b00000000000000aefffffffffffff50003e9771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc4771c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f35f11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd17c81c",
    x"070a00000000000000aefffffffffffff8ef35f2121c",
    x"080200000000000000aefffffffffffff6f669de5c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ca8f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbebd21c",
    x"020900000000000001a400000000000000fb3367611c",
    x"030b00000000000001a4fffffffffffff50003e9781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc4751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f35ee1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd17c21c",
    x"070a00000000000001a4fffffffffffff8ef35f20f1c",
    x"080200000000000001a4fffffffffffff6f669de591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ca8b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbebd31c",
    x"0209000000000000016a00000000000000fb33675b1c",
    x"030b000000000000016afffffffffffff50003e9791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc4721c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f35ea1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd17bc1c",
    x"070a000000000000016afffffffffffff8ef35f20b1c",
    x"0802000000000000016afffffffffffff6f669de571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ca861c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbebd41c",
    x"0209000000000000015500000000000000fb3367551c",
    x"030b0000000000000155fffffffffffff50003e9791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35e61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd17b61c",
    x"070a0000000000000155fffffffffffff8ef35f2071c",
    x"08020000000000000155fffffffffffff6f669de541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266ca821c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbebd51c",
    x"0209000000000000019500000000000000fb3367501c",
    x"030b0000000000000195fffffffffffff50003e97a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dc46d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f35e31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd17af1c",
    x"070a0000000000000195fffffffffffff8ef35f2031c",
    x"080200000000000002a5fffffffffffff6f669de521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ca7e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbebd61c",
    x"020900000000000002aa00000000000000fb33674a1c",
    x"030b00000000000002aafffffffffffff50003e97b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc46b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f35df1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd17a91c",
    x"070a00000000000002aafffffffffffff8ef35f2001c",
    x"08020000000000000155fffffffffffff6f669de501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266ca7a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbebd81c",
    x"0209000000000000029600000000000000fb3367441c",
    x"030b00000000000001aafffffffffffff50003e97c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc4681c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f35dc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd17a31c",
    x"070a0000000000000256fffffffffffff8ef35f1fc1c",
    x"08020000000000000155fffffffffffff6f669de4d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266ca761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbebd91c",
    x"0209000000000000026500000000000000fb33673f1c",
    x"030b00000000000002a9fffffffffffff50003e97d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc4661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f35d81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd179d1c",
    x"070a000000000000029afffffffffffff8ef35f1f81c",
    x"08020000000000000159fffffffffffff6f669de4b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266ca721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbebda1c",
    x"0209000000000000029600000000000000fb3367391c",
    x"030b000000000000016afffffffffffff50003e97e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc4631c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f35d41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd17971c",
    x"070a0000000000000159fffffffffffff8ef35f1f51c",
    x"0802000000000000015afffffffffffff6f669de481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266ca6d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbebdb1c",
    x"0209000000000000016900000000000000fb3367341c",
    x"030b0000000000000295fffffffffffff50003e97f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc4611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f35d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd17901c",
    x"070a0000000000000196fffffffffffff8ef35f1f11c",
    x"08020000000000000299fffffffffffff6f669de461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ca691c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbebdc1c",
    x"020900000000000002a500000000000000fb33672e1c",
    x"030b0000000000000156fffffffffffff50003e9801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc45e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f35cd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd178a1c",
    x"070a00000000000002a6fffffffffffff8ef35f1ed1c",
    x"080200000000000001a5fffffffffffff6f669de431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266ca651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbebdd1c",
    x"0209000000000000025500000000000000fb3367281c",
    x"030b000000000000016afffffffffffff50003e9811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc45c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f35c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd17841c",
    x"070a0000000000000295fffffffffffff8ef35f1ea1c",
    x"0802000000000000026afffffffffffff6f669de411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266ca611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbebde1c",
    x"0209000000000000029a00000000000000fb3367231c",
    x"030b0000000000000269fffffffffffff50003e9821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc4591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f35c61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd177e1c",
    x"070a0000000000000196fffffffffffff8ef35f1e61c",
    x"08020000000000000165fffffffffffff6f669de3f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266ca5d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbebdf1c",
    x"020900000000000001a600000000000000fb33671d1c",
    x"030b000000000000019afffffffffffff50003e9831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc4571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f35c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd17781c",
    x"070a000000000000026afffffffffffff8ef35f1e21c",
    x"0802000000000000019afffffffffffff6f669de3c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266ca591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbebe11c",
    x"0209000000000000025a00000000000000fb3367181c",
    x"030b00000000000002a9fffffffffffff50003e9831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc4541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f35bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd17721c",
    x"070a00000000000002a6fffffffffffff8ef35f1de1c",
    x"08020000000000000295fffffffffffff6f669de3a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266ca541c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbebe21c",
    x"0209000000000000029600000000000000fb3367121c",
    x"030b000000000000025afffffffffffff50003e9841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc4521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f35bb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd176b1c",
    x"070a000000000000019afffffffffffff8ef35f1db1c",
    x"0802000000000000029afffffffffffff6f669de371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266ca501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbebe31c",
    x"0209000000000000019900000000000000fb33670c1c",
    x"030b0000000000000156fffffffffffff50003e9851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc44f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f35b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd17651c",
    x"070a0000000000000166fffffffffffff8ef35f1d71c",
    x"080200000000000001a9fffffffffffff6f669de351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ca4c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbebe41c",
    x"0209000000000000015600000000000000fb3367071c",
    x"030b0000000000000169fffffffffffff50003e9861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc44d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f35b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd175f1c",
    x"070a0000000000000159fffffffffffff8ef35f1d31c",
    x"08020000000000000255fffffffffffff6f669de331c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266ca481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbebe51c",
    x"0209000000000000029a00000000000000fb3367011c",
    x"030b00000000000002a9fffffffffffff50003e9871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc44a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd17591c",
    x"070a0000000000000159fffffffffffff8ef35f1d01c",
    x"08020000000000000299fffffffffffff6f669de301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266ca441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbebe61c",
    x"0209000000000000031f00000000000000fb3366fb1c",
    x"030b000000000000031ffffffffffffff50003e9881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc4481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f35ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd17531c",
    x"070a000000000000031ffffffffffffff8ef35f1cc1c",
    x"0802000000000000031ffffffffffffff6f669de2e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266ca401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbebe71c",
    x"020900000000000000ae00000000000000fb3366f61c",
    x"030b00000000000000aefffffffffffff50003e9891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc4451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f35a91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd174d1c",
    x"070a00000000000000aefffffffffffff8ef35f1c81c",
    x"080200000000000000aefffffffffffff6f669de2b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266ca3b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbebe91c",
    x"020900000000000001a400000000000000fb3366f01c",
    x"030b00000000000001a4fffffffffffff50003e98a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc4431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f35a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd17461c",
    x"070a00000000000001a4fffffffffffff8ef35f1c51c",
    x"080200000000000001a4fffffffffffff6f669de291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266ca371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbebea1c",
    x"0209000000000000026a00000000000000fb3366eb1c",
    x"030b000000000000026afffffffffffff50003e98b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc4401c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f35a21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026a0000000000000004cd17401c",
    x"070a000000000000026afffffffffffff8ef35f1c11c",
    x"0802000000000000026afffffffffffff6f669de271c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ca331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbebeb1c",
    x"0209000000000000015500000000000000fb3366e51c",
    x"030b0000000000000155fffffffffffff50003e98c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc43e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f359e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd173a1c",
    x"070a00000000000002a9fffffffffffff8ef35f1bd1c",
    x"08020000000000000155fffffffffffff6f669de241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266ca2f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbebec1c",
    x"0209000000000000015500000000000000fb3366df1c",
    x"030b0000000000000155fffffffffffff50003e98d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc43b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f359a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd17341c",
    x"070a00000000000001aafffffffffffff8ef35f1b91c",
    x"08020000000000000155fffffffffffff6f669de221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266ca2b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbebed1c",
    x"0209000000000000015600000000000000fb3366da1c",
    x"030b0000000000000155fffffffffffff50003e98d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc4391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f35971c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd172e1c",
    x"070a00000000000002aafffffffffffff8ef35f1b61c",
    x"08020000000000000155fffffffffffff6f669de1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ca271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbebee1c",
    x"0209000000000000025500000000000000fb3366d41c",
    x"030b0000000000000195fffffffffffff50003e98e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc4361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f35931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd17271c",
    x"070a000000000000026afffffffffffff8ef35f1b21c",
    x"08020000000000000195fffffffffffff6f669de1d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266ca221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbebef1c",
    x"0209000000000000016500000000000000fb3366cf1c",
    x"030b00000000000002a9fffffffffffff50003e98f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc4341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35901c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002590000000000000004cd17211c",
    x"070a0000000000000256fffffffffffff8ef35f1ae1c",
    x"08020000000000000299fffffffffffff6f669de1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266ca1e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbebf01c",
    x"0209000000000000019900000000000000fb3366c91c",
    x"030b0000000000000195fffffffffffff50003e9901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc4311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f358c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd171b1c",
    x"070a0000000000000266fffffffffffff8ef35f1ab1c",
    x"080200000000000002a6fffffffffffff6f669de181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266ca1a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbebf21c",
    x"0209000000000000016500000000000000fb3366c31c",
    x"030b0000000000000166fffffffffffff50003e9911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc42f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f35881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd17151c",
    x"070a0000000000000156fffffffffffff8ef35f1a71c",
    x"0802000000000000025afffffffffffff6f669de161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266ca161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbebf31c",
    x"0209000000000000019500000000000000fb3366be1c",
    x"030b0000000000000265fffffffffffff50003e9921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc42c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f35851c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd170f1c",
    x"070a000000000000025afffffffffffff8ef35f1a31c",
    x"0802000000000000016afffffffffffff6f669de131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266ca121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbebf41c",
    x"0209000000000000026a00000000000000fb3366b81c",
    x"030b00000000000002aafffffffffffff50003e9931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc42a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f35811c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd17091c",
    x"070a0000000000000195fffffffffffff8ef35f19f1c",
    x"08020000000000000195fffffffffffff6f669de111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266ca0e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbebf51c",
    x"0209000000000000025600000000000000fb3366b21c",
    x"030b00000000000002a5fffffffffffff50003e9941c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dc4271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f357d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd17021c",
    x"070a00000000000002a5fffffffffffff8ef35f19c1c",
    x"08020000000000000295fffffffffffff6f669de0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266ca091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbebf61c",
    x"020900000000000001a900000000000000fb3366ad1c",
    x"030b0000000000000155fffffffffffff50003e9951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc4251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f357a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd16fc1c",
    x"070a0000000000000256fffffffffffff8ef35f1981c",
    x"08020000000000000199fffffffffffff6f669de0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266ca051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbebf71c",
    x"0209000000000000029500000000000000fb3366a71c",
    x"030b0000000000000299fffffffffffff50003e9961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f35761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd16f61c",
    x"070a0000000000000266fffffffffffff8ef35f1941c",
    x"08020000000000000166fffffffffffff6f669de0a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266ca011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbebf81c",
    x"0209000000000000016900000000000000fb3366a21c",
    x"030b000000000000016afffffffffffff50003e9961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc4201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f35731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd16f01c",
    x"070a0000000000000256fffffffffffff8ef35f1911c",
    x"08020000000000000199fffffffffffff6f669de071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266c9fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbebf91c",
    x"0209000000000000026a00000000000000fb33669c1c",
    x"030b000000000000016afffffffffffff50003e9971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc41d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f356f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd16ea1c",
    x"070a00000000000001a5fffffffffffff8ef35f18d1c",
    x"08020000000000000266fffffffffffff6f669de051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c9f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbebfb1c",
    x"020900000000000001a900000000000000fb3366961c",
    x"030b000000000000026afffffffffffff50003e9981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc41b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f356b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd16e41c",
    x"070a0000000000000166fffffffffffff8ef35f1891c",
    x"08020000000000000296fffffffffffff6f669de021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266c9f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbebfc1c",
    x"020900000000000002a600000000000000fb3366911c",
    x"030b000000000000015afffffffffffff50003e9991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc4181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f35681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002990000000000000004cd16dd1c",
    x"070a0000000000000295fffffffffffff8ef35f1861c",
    x"080200000000000002a5fffffffffffff6f669de001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c9f01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbebfd1c",
    x"0209000000000000031f00000000000000fb33668b1c",
    x"030b000000000000031ffffffffffffff50003e99a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc4161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f35641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd16d71c",
    x"070a000000000000031ffffffffffffff8ef35f1821c",
    x"0802000000000000031ffffffffffffff6f669ddfd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c9ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbebfe1c",
    x"020900000000000000ae00000000000000fb3366861c",
    x"030b00000000000000aefffffffffffff50003e99b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc4131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f35611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd16d11c",
    x"070a00000000000000aefffffffffffff8ef35f17e1c",
    x"080200000000000000aefffffffffffff6f669ddfb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c9e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbebff1c",
    x"020900000000000001a400000000000000fb3366801c",
    x"030b00000000000001a4fffffffffffff50003e99c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc4111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f355d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd16cb1c",
    x"070a00000000000001a4fffffffffffff8ef35f17a1c",
    x"080200000000000001a4fffffffffffff6f669ddf91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266c9e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbec001c",
    x"0209000000000000015a00000000000000fb33667a1c",
    x"030b000000000000015afffffffffffff50003e99d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc40e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f35591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd16c51c",
    x"070a000000000000015afffffffffffff8ef35f1771c",
    x"0802000000000000015afffffffffffff6f669ddf61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec011c",
    x"020900000000000001aa00000000000000fb3366751c",
    x"030b0000000000000255fffffffffffff50003e99e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc40c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd16be1c",
    x"070a0000000000000155fffffffffffff8ef35f1731c",
    x"08020000000000000155fffffffffffff6f669ddf41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266c9dc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbec031c",
    x"0209000000000000016900000000000000fb33666f1c",
    x"030b0000000000000269fffffffffffff50003e99f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc4091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f35521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd16b81c",
    x"070a00000000000002a6fffffffffffff8ef35f16f1c",
    x"080200000000000001a5fffffffffffff6f669ddf11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266c9d71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbec041c",
    x"020900000000000001a600000000000000fb3366691c",
    x"030b0000000000000296fffffffffffff50003e9a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc4071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f354e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd16b21c",
    x"070a000000000000029afffffffffffff8ef35f16c1c",
    x"08020000000000000196fffffffffffff6f669ddef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c9d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbec051c",
    x"0209000000000000026900000000000000fb3366641c",
    x"030b0000000000000255fffffffffffff50003e9a01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc4041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f354b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001990000000000000004cd16ac1c",
    x"070a0000000000000265fffffffffffff8ef35f1681c",
    x"08020000000000000256fffffffffffff6f669dded1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbec061c",
    x"0209000000000000015600000000000000fb33665e1c",
    x"030b0000000000000155fffffffffffff50003e9a11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc4021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f35471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd16a61c",
    x"070a00000000000002aafffffffffffff8ef35f1641c",
    x"08020000000000000155fffffffffffff6f669ddea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266c9cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbec071c",
    x"0209000000000000026500000000000000fb3366591c",
    x"030b0000000000000265fffffffffffff50003e9a21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc3ff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f35441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002650000000000000004cd16a01c",
    x"070a000000000000019afffffffffffff8ef35f1601c",
    x"08020000000000000265fffffffffffff6f669dde81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec081c",
    x"020900000000000002aa00000000000000fb3366531c",
    x"030b00000000000002aafffffffffffff50003e9a31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3fd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16991c",
    x"070a0000000000000155fffffffffffff8ef35f15d1c",
    x"080200000000000002aafffffffffffff6f669dde51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec091c",
    x"020900000000000002aa00000000000000fb33664d1c",
    x"030b00000000000002aafffffffffffff50003e9a41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3fa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f353c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16931c",
    x"070a0000000000000155fffffffffffff8ef35f1591c",
    x"080200000000000002aafffffffffffff6f669dde31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec0a1c",
    x"020900000000000002aa00000000000000fb3366481c",
    x"030b00000000000002aafffffffffffff50003e9a51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd168d1c",
    x"070a0000000000000155fffffffffffff8ef35f1551c",
    x"080200000000000002aafffffffffffff6f669dde11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266c9ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbec0c1c",
    x"020900000000000001a600000000000000fb3366421c",
    x"030b00000000000001a6fffffffffffff50003e9a61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000259fffffffffffff4099dc3f51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f35351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd16871c",
    x"070a0000000000000259fffffffffffff8ef35f1521c",
    x"080200000000000001a6fffffffffffff6f669ddde1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec0d1c",
    x"020900000000000002aa00000000000000fb33663d1c",
    x"030b00000000000002aafffffffffffff50003e9a71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3f31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f35321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16811c",
    x"070a0000000000000155fffffffffffff8ef35f14e1c",
    x"080200000000000002aafffffffffffff6f669dddc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec0e1c",
    x"020900000000000002aa00000000000000fb3366371c",
    x"030b00000000000002aafffffffffffff50003e9a81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3f01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f352e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd167a1c",
    x"070a0000000000000155fffffffffffff8ef35f14a1c",
    x"080200000000000002aafffffffffffff6f669ddd91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c9ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbec0f1c",
    x"020900000000000002a600000000000000fb3366311c",
    x"030b00000000000002a6fffffffffffff50003e9a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc3ee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f352a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd16741c",
    x"070a0000000000000159fffffffffffff8ef35f1471c",
    x"080200000000000002a6fffffffffffff6f669ddd71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c9aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a50000000000000b0bfbec101c",
    x"0209000000000000029500000000000000fb33662c1c",
    x"030b00000000000002aafffffffffffff50003e9a91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc3eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f35271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd166e1c",
    x"070a000000000000019afffffffffffff8ef35f1431c",
    x"080200000000000002a5fffffffffffff6f669ddd41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec111c",
    x"0209000000000000026a00000000000000fb3366261c",
    x"030b000000000000026afffffffffffff50003e9aa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc3e91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f35231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002650000000000000004cd16681c",
    x"070a0000000000000165fffffffffffff8ef35f13f1c",
    x"080200000000000002aafffffffffffff6f669ddd21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266c9a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec121c",
    x"0209000000000000015600000000000000fb3366201c",
    x"030b0000000000000156fffffffffffff50003e9ab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dc3e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f351f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd16621c",
    x"070a00000000000002a9fffffffffffff8ef35f13b1c",
    x"08020000000000000156fffffffffffff6f669ddd01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c99d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec141c",
    x"0209000000000000031f00000000000000fb33661b1c",
    x"030b000000000000031ffffffffffffff50003e9ac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc3e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f351c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd165c1c",
    x"070a000000000000031ffffffffffffff8ef35f1381c",
    x"0802000000000000031ffffffffffffff6f669ddcd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c9991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec151c",
    x"020900000000000000ae00000000000000fb3366151c",
    x"030b00000000000000aefffffffffffff50003e9ad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc3e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f35181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd16551c",
    x"070a00000000000000aefffffffffffff8ef35f1341c",
    x"080200000000000000aefffffffffffff6f669ddcb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c9951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec161c",
    x"020900000000000001a400000000000000fb3366101c",
    x"030b00000000000001a4fffffffffffff50003e9ae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc3df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f35151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd164f1c",
    x"070a00000000000001a4fffffffffffff8ef35f1301c",
    x"080200000000000001a4fffffffffffff6f669ddc81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266c9911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbec171c",
    x"0209000000000000025a00000000000000fb33660a1c",
    x"030b000000000000025afffffffffffff50003e9af1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc3dc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f35111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd16491c",
    x"070a000000000000025afffffffffffff8ef35f12d1c",
    x"0802000000000000025afffffffffffff6f669ddc61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c98c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec181c",
    x"020900000000000002aa00000000000000fb3366041c",
    x"030b00000000000002aafffffffffffff50003e9b01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f350d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16431c",
    x"070a00000000000002aafffffffffffff8ef35f1291c",
    x"080200000000000002aafffffffffffff6f669ddc41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c9881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbec191c",
    x"0209000000000000029a00000000000000fb3365ff1c",
    x"030b000000000000029afffffffffffff50003e9b11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc3d71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f350a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd163d1c",
    x"070a000000000000029afffffffffffff8ef35f1251c",
    x"0802000000000000029afffffffffffff6f669ddc11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec1a1c",
    x"020900000000000002aa00000000000000fb3365f91c",
    x"030b00000000000002aafffffffffffff50003e9b21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3d51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f35061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16361c",
    x"070a00000000000002aafffffffffffff8ef35f1211c",
    x"080200000000000002aafffffffffffff6f669ddbf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec1b1c",
    x"020900000000000002aa00000000000000fb3365f41c",
    x"030b00000000000002aafffffffffffff50003e9b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3d21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f35031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16301c",
    x"070a00000000000002aafffffffffffff8ef35f11e1c",
    x"080200000000000002aafffffffffffff6f669ddbc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c97c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec1d1c",
    x"020900000000000002aa00000000000000fb3365ee1c",
    x"030b00000000000002aafffffffffffff50003e9b31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3d01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd162a1c",
    x"070a00000000000002aafffffffffffff8ef35f11a1c",
    x"080200000000000002aafffffffffffff6f669ddba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec1e1c",
    x"020900000000000002aa00000000000000fb3365e81c",
    x"030b00000000000002aafffffffffffff50003e9b41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3cd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16241c",
    x"070a00000000000002aafffffffffffff8ef35f1161c",
    x"080200000000000002aafffffffffffff6f669ddb71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec1f1c",
    x"020900000000000002aa00000000000000fb3365e31c",
    x"030b00000000000002aafffffffffffff50003e9b51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3cb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd161e1c",
    x"070a00000000000002aafffffffffffff8ef35f1131c",
    x"080200000000000002aafffffffffffff6f669ddb51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c96f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec201c",
    x"020900000000000002aa00000000000000fb3365dd1c",
    x"030b00000000000002aafffffffffffff50003e9b61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3c81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16181c",
    x"070a00000000000002aafffffffffffff8ef35f10f1c",
    x"080200000000000002aafffffffffffff6f669ddb31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c96b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec211c",
    x"020900000000000002aa00000000000000fb3365d71c",
    x"030b00000000000002aafffffffffffff50003e9b71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3c61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd16111c",
    x"070a00000000000002aafffffffffffff8ef35f10b1c",
    x"080200000000000002aafffffffffffff6f669ddb01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266c9671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbec221c",
    x"0209000000000000016600000000000000fb3365d21c",
    x"030b0000000000000166fffffffffffff50003e9b81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc3c31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f34ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd160b1c",
    x"070a0000000000000166fffffffffffff8ef35f1081c",
    x"08020000000000000166fffffffffffff6f669ddae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec231c",
    x"0209000000000000015500000000000000fb3365cc1c",
    x"030b0000000000000155fffffffffffff50003e9b91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3c11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd16051c",
    x"070a0000000000000155fffffffffffff8ef35f1041c",
    x"08020000000000000155fffffffffffff6f669ddab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c95f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec251c",
    x"0209000000000000015500000000000000fb3365c71c",
    x"030b0000000000000155fffffffffffff50003e9ba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3be1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34e61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15ff1c",
    x"070a0000000000000155fffffffffffff8ef35f1001c",
    x"08020000000000000155fffffffffffff6f669dda91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c95a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec261c",
    x"0209000000000000015500000000000000fb3365c11c",
    x"030b0000000000000155fffffffffffff50003e9bb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3bc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15f91c",
    x"070a0000000000000155fffffffffffff8ef35f0fc1c",
    x"08020000000000000155fffffffffffff6f669dda71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec271c",
    x"0209000000000000015500000000000000fb3365bb1c",
    x"030b0000000000000155fffffffffffff50003e9bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3b91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15f31c",
    x"070a0000000000000155fffffffffffff8ef35f0f91c",
    x"08020000000000000155fffffffffffff6f669dda41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c9521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec281c",
    x"0209000000000000015500000000000000fb3365b61c",
    x"030b0000000000000155fffffffffffff50003e9bc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3b71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34db1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15ec1c",
    x"070a0000000000000155fffffffffffff8ef35f0f51c",
    x"08020000000000000155fffffffffffff6f669dda21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c94e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbec291c",
    x"0209000000000000015900000000000000fb3365b01c",
    x"030b0000000000000159fffffffffffff50003e9bd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc3b41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f34d71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd15e61c",
    x"070a0000000000000159fffffffffffff8ef35f0f11c",
    x"08020000000000000159fffffffffffff6f669dd9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c94a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec2a1c",
    x"0209000000000000031f00000000000000fb3365ab1c",
    x"030b000000000000031ffffffffffffff50003e9be1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc3b21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f34d41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd15e01c",
    x"070a000000000000031ffffffffffffff8ef35f0ee1c",
    x"0802000000000000031ffffffffffffff6f669dd9d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c9461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec2b1c",
    x"020900000000000000ae00000000000000fb3365a51c",
    x"030b00000000000000aefffffffffffff50003e9bf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc3af1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f34d01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd15da1c",
    x"070a00000000000000aefffffffffffff8ef35f0ea1c",
    x"080200000000000000aefffffffffffff6f669dd9b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c9411c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec2c1c",
    x"020900000000000001a400000000000000fb33659f1c",
    x"030b00000000000001a4fffffffffffff50003e9c01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc3ad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f34cc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd15d41c",
    x"070a00000000000001a4fffffffffffff8ef35f0e61c",
    x"080200000000000001a4fffffffffffff6f669dd981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c93d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbec2e1c",
    x"0209000000000000029a00000000000000fb33659a1c",
    x"030b000000000000029afffffffffffff50003e9c11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc3aa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f34c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd15cd1c",
    x"070a000000000000029afffffffffffff8ef35f0e21c",
    x"0802000000000000029afffffffffffff6f669dd961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec2f1c",
    x"020900000000000002aa00000000000000fb3365941c",
    x"030b00000000000002aafffffffffffff50003e9c21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3a81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34c51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15c71c",
    x"070a00000000000002aafffffffffffff8ef35f0df1c",
    x"080200000000000002aafffffffffffff6f669dd931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c9351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbec301c",
    x"0209000000000000029a00000000000000fb33658e1c",
    x"030b000000000000029afffffffffffff50003e9c31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc3a51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f34c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd15c11c",
    x"070a000000000000029afffffffffffff8ef35f0db1c",
    x"0802000000000000029afffffffffffff6f669dd911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec311c",
    x"020900000000000002aa00000000000000fb3365891c",
    x"030b00000000000002aafffffffffffff50003e9c41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3a31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15bb1c",
    x"070a00000000000002aafffffffffffff8ef35f0d71c",
    x"080200000000000002aafffffffffffff6f669dd8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c92d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec321c",
    x"020900000000000002aa00000000000000fb3365831c",
    x"030b00000000000002aafffffffffffff50003e9c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3a01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34ba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15b51c",
    x"070a00000000000002aafffffffffffff8ef35f0d41c",
    x"080200000000000002aafffffffffffff6f669dd8c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9281c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec331c",
    x"020900000000000002aa00000000000000fb33657e1c",
    x"030b00000000000002aafffffffffffff50003e9c51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc39e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15af1c",
    x"070a00000000000002aafffffffffffff8ef35f0d01c",
    x"080200000000000002aafffffffffffff6f669dd8a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec341c",
    x"020900000000000002aa00000000000000fb3365781c",
    x"030b00000000000002aafffffffffffff50003e9c61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc39b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15a81c",
    x"070a00000000000002aafffffffffffff8ef35f0cc1c",
    x"080200000000000002aafffffffffffff6f669dd871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec361c",
    x"020900000000000002aa00000000000000fb3365721c",
    x"030b00000000000002aafffffffffffff50003e9c71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3991c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34af1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15a21c",
    x"070a00000000000002aafffffffffffff8ef35f0c81c",
    x"080200000000000002aafffffffffffff6f669dd851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c91c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec371c",
    x"020900000000000002aa00000000000000fb33656d1c",
    x"030b00000000000002aafffffffffffff50003e9c81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd159c1c",
    x"070a00000000000002aafffffffffffff8ef35f0c51c",
    x"080200000000000002aafffffffffffff6f669dd821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec381c",
    x"020900000000000002aa00000000000000fb3365671c",
    x"030b00000000000002aafffffffffffff50003e9c91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3941c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15961c",
    x"070a00000000000002aafffffffffffff8ef35f0c11c",
    x"080200000000000002aafffffffffffff6f669dd801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec391c",
    x"020900000000000002aa00000000000000fb3365621c",
    x"030b00000000000002aafffffffffffff50003e9ca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15901c",
    x"070a00000000000002aafffffffffffff8ef35f0bd1c",
    x"080200000000000002aafffffffffffff6f669dd7e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec3a1c",
    x"020900000000000002aa00000000000000fb33655c1c",
    x"030b00000000000002aafffffffffffff50003e9cb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc38f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15891c",
    x"070a00000000000002aafffffffffffff8ef35f0ba1c",
    x"080200000000000002aafffffffffffff6f669dd7b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c90b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec3b1c",
    x"020900000000000002aa00000000000000fb3365561c",
    x"030b00000000000002aafffffffffffff50003e9cc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc38c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f349d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15831c",
    x"070a00000000000002aafffffffffffff8ef35f0b61c",
    x"080200000000000002aafffffffffffff6f669dd791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec3c1c",
    x"020900000000000002aa00000000000000fb3365511c",
    x"030b00000000000002aafffffffffffff50003e9cd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc38a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f349a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd157d1c",
    x"070a00000000000002aafffffffffffff8ef35f0b21c",
    x"080200000000000002aafffffffffffff6f669dd761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c9031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec3d1c",
    x"020900000000000002aa00000000000000fb33654b1c",
    x"030b00000000000002aafffffffffffff50003e9ce1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f34961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd15771c",
    x"070a00000000000002aafffffffffffff8ef35f0ae1c",
    x"080200000000000002aafffffffffffff6f669dd741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266c8ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbec3f1c",
    x"020900000000000001aa00000000000000fb3365451c",
    x"030b00000000000001aafffffffffffff50003e9ce1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc3851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f34931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd15711c",
    x"070a00000000000001aafffffffffffff8ef35f0ab1c",
    x"080200000000000001aafffffffffffff6f669dd711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8fb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec401c",
    x"0209000000000000015500000000000000fb3365401c",
    x"030b0000000000000155fffffffffffff50003e9cf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f348f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd156b1c",
    x"070a0000000000000155fffffffffffff8ef35f0a71c",
    x"08020000000000000155fffffffffffff6f669dd6f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c8f71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec411c",
    x"0209000000000000031f00000000000000fb33653a1c",
    x"030b000000000000031ffffffffffffff50003e9d01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc3801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f348b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd15641c",
    x"070a000000000000031ffffffffffffff8ef35f0a31c",
    x"0802000000000000031ffffffffffffff6f669dd6d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c8f21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec421c",
    x"020900000000000000ae00000000000000fb3365351c",
    x"030b00000000000000aefffffffffffff50003e9d11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc37d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f34881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd155e1c",
    x"070a00000000000000aefffffffffffff8ef35f0a01c",
    x"080200000000000000aefffffffffffff6f669dd6a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c8ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec431c",
    x"020900000000000001a400000000000000fb33652f1c",
    x"030b00000000000001a4fffffffffffff50003e9d21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc37b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f34841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd15581c",
    x"070a00000000000001a4fffffffffffff8ef35f09c1c",
    x"080200000000000001a4fffffffffffff6f669dd681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266c8ea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbec441c",
    x"0209000000000000019a00000000000000fb3365291c",
    x"030b000000000000019afffffffffffff50003e9d31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc3781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f34811c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd15521c",
    x"070a000000000000019afffffffffffff8ef35f0981c",
    x"0802000000000000019afffffffffffff6f669dd651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8e61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec451c",
    x"0209000000000000015500000000000000fb3365241c",
    x"030b0000000000000155fffffffffffff50003e9d41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f347d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd154c1c",
    x"070a0000000000000155fffffffffffff8ef35f0941c",
    x"08020000000000000155fffffffffffff6f669dd631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8e21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec471c",
    x"0209000000000000015500000000000000fb33651e1c",
    x"030b0000000000000155fffffffffffff50003e9d51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15451c",
    x"070a0000000000000155fffffffffffff8ef35f0911c",
    x"08020000000000000155fffffffffffff6f669dd611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8de1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec481c",
    x"0209000000000000015500000000000000fb3365191c",
    x"030b0000000000000155fffffffffffff50003e9d61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd153f1c",
    x"070a0000000000000155fffffffffffff8ef35f08d1c",
    x"08020000000000000155fffffffffffff6f669dd5e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8d91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec491c",
    x"0209000000000000015500000000000000fb3365131c",
    x"030b0000000000000155fffffffffffff50003e9d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc36e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15391c",
    x"070a0000000000000155fffffffffffff8ef35f0891c",
    x"08020000000000000155fffffffffffff6f669dd5c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8d51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec4a1c",
    x"0209000000000000015500000000000000fb33650d1c",
    x"030b0000000000000155fffffffffffff50003e9d71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc36c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f346e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15331c",
    x"070a0000000000000155fffffffffffff8ef35f0861c",
    x"08020000000000000155fffffffffffff6f669dd591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8d11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec4b1c",
    x"0209000000000000015500000000000000fb3365081c",
    x"030b0000000000000155fffffffffffff50003e9d81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f346b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd152d1c",
    x"070a0000000000000155fffffffffffff8ef35f0821c",
    x"08020000000000000155fffffffffffff6f669dd571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8cd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec4c1c",
    x"0209000000000000015500000000000000fb3365021c",
    x"030b0000000000000155fffffffffffff50003e9d91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15271c",
    x"070a0000000000000155fffffffffffff8ef35f07e1c",
    x"08020000000000000155fffffffffffff6f669dd541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8c91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec4d1c",
    x"0209000000000000015500000000000000fb3364fc1c",
    x"030b0000000000000155fffffffffffff50003e9da1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15201c",
    x"070a0000000000000155fffffffffffff8ef35f07b1c",
    x"08020000000000000155fffffffffffff6f669dd521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8c51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec4f1c",
    x"0209000000000000015500000000000000fb3364f71c",
    x"030b0000000000000155fffffffffffff50003e9db1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34601c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd151a1c",
    x"070a0000000000000155fffffffffffff8ef35f0771c",
    x"08020000000000000155fffffffffffff6f669dd501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8c01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec501c",
    x"0209000000000000015500000000000000fb3364f11c",
    x"030b0000000000000155fffffffffffff50003e9dc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc35f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f345c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15141c",
    x"070a0000000000000155fffffffffffff8ef35f0731c",
    x"08020000000000000155fffffffffffff6f669dd4d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8bc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec511c",
    x"0209000000000000015500000000000000fb3364ec1c",
    x"030b0000000000000155fffffffffffff50003e9dd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc35c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd150e1c",
    x"070a0000000000000155fffffffffffff8ef35f06f1c",
    x"08020000000000000155fffffffffffff6f669dd4b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8b81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec521c",
    x"0209000000000000015500000000000000fb3364e61c",
    x"030b0000000000000155fffffffffffff50003e9de1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc35a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15081c",
    x"070a0000000000000155fffffffffffff8ef35f06c1c",
    x"08020000000000000155fffffffffffff6f669dd481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8b41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec531c",
    x"0209000000000000015500000000000000fb3364e01c",
    x"030b0000000000000155fffffffffffff50003e9df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd15011c",
    x"070a0000000000000155fffffffffffff8ef35f0681c",
    x"08020000000000000155fffffffffffff6f669dd461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8b01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec541c",
    x"0209000000000000015500000000000000fb3364db1c",
    x"030b0000000000000155fffffffffffff50003e9df1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f344e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14fb1c",
    x"070a0000000000000155fffffffffffff8ef35f0641c",
    x"08020000000000000155fffffffffffff6f669dd441c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8ac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec551c",
    x"0209000000000000015500000000000000fb3364d51c",
    x"030b0000000000000155fffffffffffff50003e9e01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f344a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14f51c",
    x"070a0000000000000155fffffffffffff8ef35f0611c",
    x"08020000000000000155fffffffffffff6f669dd411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8a71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec561c",
    x"0209000000000000015500000000000000fb3364cf1c",
    x"030b0000000000000155fffffffffffff50003e9e11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14ef1c",
    x"070a0000000000000155fffffffffffff8ef35f05d1c",
    x"08020000000000000155fffffffffffff6f669dd3f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c8a31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec581c",
    x"0209000000000000031f00000000000000fb3364ca1c",
    x"030b000000000000031ffffffffffffff50003e9e21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc34d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f34431c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd14e91c",
    x"070a000000000000031ffffffffffffff8ef35f0591c",
    x"0802000000000000031ffffffffffffff6f669dd3c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c89f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec591c",
    x"020900000000000000ae00000000000000fb3364c41c",
    x"030b00000000000000aefffffffffffff50003e9e31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc34b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f34401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd14e31c",
    x"070a00000000000000aefffffffffffff8ef35f0551c",
    x"080200000000000000aefffffffffffff6f669dd3a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c89b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec5a1c",
    x"020900000000000001a400000000000000fb3364bf1c",
    x"030b00000000000001a4fffffffffffff50003e9e41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc3481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f343c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd14dc1c",
    x"070a00000000000001a4fffffffffffff8ef35f0521c",
    x"080200000000000001a4fffffffffffff6f669dd371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266c8971c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbec5b1c",
    x"0209000000000000015600000000000000fb3364b91c",
    x"030b0000000000000156fffffffffffff50003e9e51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc3461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f34381c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd14d61c",
    x"070a0000000000000156fffffffffffff8ef35f04e1c",
    x"08020000000000000156fffffffffffff6f669dd351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c8931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbec5c1c",
    x"0209000000000000029500000000000000fb3364b31c",
    x"030b0000000000000295fffffffffffff50003e9e61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc3431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f34351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd14d01c",
    x"070a0000000000000295fffffffffffff8ef35f04a1c",
    x"08020000000000000295fffffffffffff6f669dd331c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c88e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec5d1c",
    x"0209000000000000015500000000000000fb3364ae1c",
    x"030b0000000000000155fffffffffffff50003e9e71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34311c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14ca1c",
    x"070a0000000000000155fffffffffffff8ef35f0471c",
    x"08020000000000000155fffffffffffff6f669dd301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c88a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec5e1c",
    x"0209000000000000015500000000000000fb3364a81c",
    x"030b0000000000000155fffffffffffff50003e9e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc33e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f342e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14c41c",
    x"070a0000000000000155fffffffffffff8ef35f0431c",
    x"08020000000000000155fffffffffffff6f669dd2e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8861c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec601c",
    x"0209000000000000015500000000000000fb3364a31c",
    x"030b0000000000000155fffffffffffff50003e9e81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc33c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f342a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14bd1c",
    x"070a0000000000000155fffffffffffff8ef35f03f1c",
    x"08020000000000000155fffffffffffff6f669dd2b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8821c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec611c",
    x"0209000000000000015500000000000000fb33649d1c",
    x"030b0000000000000155fffffffffffff50003e9e91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34261c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14b71c",
    x"070a0000000000000155fffffffffffff8ef35f03b1c",
    x"08020000000000000155fffffffffffff6f669dd291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c87e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec621c",
    x"0209000000000000015500000000000000fb3364971c",
    x"030b0000000000000155fffffffffffff50003e9ea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14b11c",
    x"070a0000000000000155fffffffffffff8ef35f0381c",
    x"08020000000000000155fffffffffffff6f669dd271c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c87a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec631c",
    x"0209000000000000015500000000000000fb3364921c",
    x"030b0000000000000155fffffffffffff50003e9eb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f341f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14ab1c",
    x"070a0000000000000155fffffffffffff8ef35f0341c",
    x"08020000000000000155fffffffffffff6f669dd241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8751c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec641c",
    x"0209000000000000015500000000000000fb33648c1c",
    x"030b0000000000000155fffffffffffff50003e9ec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f341b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14a51c",
    x"070a0000000000000155fffffffffffff8ef35f0301c",
    x"08020000000000000155fffffffffffff6f669dd221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8711c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec651c",
    x"0209000000000000015500000000000000fb3364861c",
    x"030b0000000000000155fffffffffffff50003e9ed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc32f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd149f1c",
    x"070a0000000000000155fffffffffffff8ef35f02d1c",
    x"08020000000000000155fffffffffffff6f669dd1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c86d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec661c",
    x"0209000000000000015500000000000000fb3364811c",
    x"030b0000000000000155fffffffffffff50003e9ee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc32d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14981c",
    x"070a0000000000000155fffffffffffff8ef35f0291c",
    x"08020000000000000155fffffffffffff6f669dd1d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8691c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec671c",
    x"0209000000000000015500000000000000fb33647b1c",
    x"030b0000000000000155fffffffffffff50003e9ef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc32a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14921c",
    x"070a0000000000000155fffffffffffff8ef35f0251c",
    x"08020000000000000155fffffffffffff6f669dd1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec691c",
    x"0209000000000000015500000000000000fb3364761c",
    x"030b0000000000000155fffffffffffff50003e9f01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f340d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd148c1c",
    x"070a0000000000000155fffffffffffff8ef35f0211c",
    x"08020000000000000155fffffffffffff6f669dd181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c8611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec6a1c",
    x"0209000000000000015500000000000000fb3364701c",
    x"030b0000000000000155fffffffffffff50003e9f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14861c",
    x"070a0000000000000155fffffffffffff8ef35f01e1c",
    x"08020000000000000155fffffffffffff6f669dd161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c85d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec6b1c",
    x"0209000000000000015500000000000000fb33646a1c",
    x"030b0000000000000155fffffffffffff50003e9f11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc3231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f34061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd14801c",
    x"070a0000000000000155fffffffffffff8ef35f01a1c",
    x"08020000000000000155fffffffffffff6f669dd131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266c8581c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbec6c1c",
    x"0209000000000000019500000000000000fb3364651c",
    x"030b0000000000000195fffffffffffff50003e9f21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dc3201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f34021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001950000000000000004cd14791c",
    x"070a0000000000000195fffffffffffff8ef35f0161c",
    x"08020000000000000195fffffffffffff6f669dd111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8541c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec6d1c",
    x"020900000000000002aa00000000000000fb33645f1c",
    x"030b00000000000002aafffffffffffff50003e9f31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc31e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14731c",
    x"070a00000000000002aafffffffffffff8ef35f0131c",
    x"080200000000000002aafffffffffffff6f669dd0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c8501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec6e1c",
    x"0209000000000000031f00000000000000fb33645a1c",
    x"030b000000000000031ffffffffffffff50003e9f41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc31b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f33fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd146d1c",
    x"070a000000000000031ffffffffffffff8ef35f00f1c",
    x"0802000000000000031ffffffffffffff6f669dd0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c84c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec6f1c",
    x"020900000000000000ae00000000000000fb3364541c",
    x"030b00000000000000aefffffffffffff50003e9f51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc3191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f33f71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd14671c",
    x"070a00000000000000aefffffffffffff8ef35f00b1c",
    x"080200000000000000aefffffffffffff6f669dd0a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c8481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec711c",
    x"020900000000000001a400000000000000fb33644e1c",
    x"030b00000000000001a4fffffffffffff50003e9f61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc3161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f33f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd14611c",
    x"070a00000000000001a4fffffffffffff8ef35f0071c",
    x"080200000000000001a4fffffffffffff6f669dd071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266c8441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbec721c",
    x"0209000000000000025600000000000000fb3364491c",
    x"030b0000000000000256fffffffffffff50003e9f71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dc3141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f33f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd145b1c",
    x"070a0000000000000256fffffffffffff8ef35f0041c",
    x"08020000000000000256fffffffffffff6f669dd051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c83f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec731c",
    x"020900000000000002aa00000000000000fb3364431c",
    x"030b00000000000002aafffffffffffff50003e9f81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14541c",
    x"070a00000000000002aafffffffffffff8ef35f0001c",
    x"080200000000000002aafffffffffffff6f669dd021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c83b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec741c",
    x"020900000000000002aa00000000000000fb33643d1c",
    x"030b00000000000002aafffffffffffff50003e9f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc30f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd144e1c",
    x"070a00000000000002aafffffffffffff8ef35effc1c",
    x"080200000000000002aafffffffffffff6f669dd001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec751c",
    x"020900000000000002aa00000000000000fb3364381c",
    x"030b00000000000002aafffffffffffff50003e9f91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc30c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33e51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14481c",
    x"070a00000000000002aafffffffffffff8ef35eff81c",
    x"080200000000000002aafffffffffffff6f669dcfd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec761c",
    x"020900000000000002aa00000000000000fb3364321c",
    x"030b00000000000002aafffffffffffff50003e9fa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc30a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14421c",
    x"070a00000000000002aafffffffffffff8ef35eff51c",
    x"080200000000000002aafffffffffffff6f669dcfb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c82f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec771c",
    x"020900000000000002aa00000000000000fb33642d1c",
    x"030b00000000000002aafffffffffffff50003e9fb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd143c1c",
    x"070a00000000000002aafffffffffffff8ef35eff11c",
    x"080200000000000002aafffffffffffff6f669dcf91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c82b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec791c",
    x"020900000000000002aa00000000000000fb3364271c",
    x"030b00000000000002aafffffffffffff50003e9fc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33db1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14351c",
    x"070a00000000000002aafffffffffffff8ef35efed1c",
    x"080200000000000002aafffffffffffff6f669dcf61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec7a1c",
    x"020900000000000002aa00000000000000fb3364211c",
    x"030b00000000000002aafffffffffffff50003e9fd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33d71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd142f1c",
    x"070a00000000000002aafffffffffffff8ef35efea1c",
    x"080200000000000002aafffffffffffff6f669dcf41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec7b1c",
    x"020900000000000002aa00000000000000fb33641c1c",
    x"030b00000000000002aafffffffffffff50003e9fe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc3001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33d31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14291c",
    x"070a00000000000002aafffffffffffff8ef35efe61c",
    x"080200000000000002aafffffffffffff6f669dcf11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c81e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec7c1c",
    x"020900000000000002aa00000000000000fb3364161c",
    x"030b00000000000002aafffffffffffff50003e9ff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2fd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33d01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14231c",
    x"070a00000000000002aafffffffffffff8ef35efe21c",
    x"080200000000000002aafffffffffffff6f669dcef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c81a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec7d1c",
    x"020900000000000002aa00000000000000fb3364111c",
    x"030b00000000000002aafffffffffffff50003ea001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2fb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33cc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd141d1c",
    x"070a00000000000002aafffffffffffff8ef35efde1c",
    x"080200000000000002aafffffffffffff6f669dced1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec7e1c",
    x"020900000000000002aa00000000000000fb33640b1c",
    x"030b00000000000002aafffffffffffff50003ea011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33c81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14171c",
    x"070a00000000000002aafffffffffffff8ef35efdb1c",
    x"080200000000000002aafffffffffffff6f669dcea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec7f1c",
    x"020900000000000002aa00000000000000fb3364051c",
    x"030b00000000000002aafffffffffffff50003ea011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2f61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33c51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14101c",
    x"070a00000000000002aafffffffffffff8ef35efd71c",
    x"080200000000000002aafffffffffffff6f669dce81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c80d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec801c",
    x"020900000000000002aa00000000000000fb3364001c",
    x"030b00000000000002aafffffffffffff50003ea021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2f31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33c11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd140a1c",
    x"070a00000000000002aafffffffffffff8ef35efd31c",
    x"080200000000000002aafffffffffffff6f669dce51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec821c",
    x"020900000000000002aa00000000000000fb3363fa1c",
    x"030b00000000000002aafffffffffffff50003ea031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2f11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd14041c",
    x"070a00000000000002aafffffffffffff8ef35efd01c",
    x"080200000000000002aafffffffffffff6f669dce31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c8051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbec831c",
    x"0209000000000000029a00000000000000fb3363f41c",
    x"030b000000000000029afffffffffffff50003ea041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc2ee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f33ba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd13fe1c",
    x"070a000000000000029afffffffffffff8ef35efcc1c",
    x"0802000000000000029afffffffffffff6f669dce01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c8011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec841c",
    x"020900000000000002aa00000000000000fb3363ef1c",
    x"030b00000000000002aafffffffffffff50003ea051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33b61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd13f81c",
    x"070a00000000000002aafffffffffffff8ef35efc81c",
    x"080200000000000002aafffffffffffff6f669dcde1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c7fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec851c",
    x"0209000000000000031f00000000000000fb3363e91c",
    x"030b000000000000031ffffffffffffff50003ea061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc2e91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f33b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd13f11c",
    x"070a000000000000031ffffffffffffff8ef35efc41c",
    x"0802000000000000031ffffffffffffff6f669dcdc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c7f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec861c",
    x"020900000000000000ae00000000000000fb3363e41c",
    x"030b00000000000000aefffffffffffff50003ea071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc2e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f33af1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd13eb1c",
    x"070a00000000000000aefffffffffffff8ef35efc11c",
    x"080200000000000000aefffffffffffff6f669dcd91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c7f41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec871c",
    x"020900000000000001a400000000000000fb3363de1c",
    x"030b00000000000001a4fffffffffffff50003ea081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc2e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f33ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd13e51c",
    x"070a00000000000001a4fffffffffffff8ef35efbd1c",
    x"080200000000000001a4fffffffffffff6f669dcd71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266c7f01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbec881c",
    x"0209000000000000029600000000000000fb3363d81c",
    x"030b0000000000000296fffffffffffff50003ea091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dc2e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f33a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd13df1c",
    x"070a0000000000000296fffffffffffff8ef35efb91c",
    x"08020000000000000296fffffffffffff6f669dcd41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c7ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbec8a1c",
    x"020900000000000002aa00000000000000fb3363d31c",
    x"030b00000000000002aafffffffffffff50003ea0a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2df1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33a41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd13d91c",
    x"070a00000000000002aafffffffffffff8ef35efb61c",
    x"080200000000000002aafffffffffffff6f669dcd21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266c7e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbec8b1c",
    x"0209000000000000016500000000000000fb3363cd1c",
    x"030b0000000000000165fffffffffffff50003ea0a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc2dc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f33a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd13d31c",
    x"070a0000000000000165fffffffffffff8ef35efb21c",
    x"08020000000000000165fffffffffffff6f669dcd01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec8c1c",
    x"0209000000000000015500000000000000fb3363c71c",
    x"030b0000000000000155fffffffffffff50003ea0b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2da1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f339d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13cc1c",
    x"070a0000000000000155fffffffffffff8ef35efae1c",
    x"08020000000000000155fffffffffffff6f669dccd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec8d1c",
    x"0209000000000000015500000000000000fb3363c21c",
    x"030b0000000000000155fffffffffffff50003ea0c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2d71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f339a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13c61c",
    x"070a0000000000000155fffffffffffff8ef35efaa1c",
    x"08020000000000000155fffffffffffff6f669dccb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7db1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec8e1c",
    x"0209000000000000015500000000000000fb3363bc1c",
    x"030b0000000000000155fffffffffffff50003ea0d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2d51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13c01c",
    x"070a0000000000000155fffffffffffff8ef35efa71c",
    x"08020000000000000155fffffffffffff6f669dcc81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7d71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec8f1c",
    x"0209000000000000015500000000000000fb3363b71c",
    x"030b0000000000000155fffffffffffff50003ea0e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2d21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13ba1c",
    x"070a0000000000000155fffffffffffff8ef35efa31c",
    x"08020000000000000155fffffffffffff6f669dcc61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec901c",
    x"0209000000000000015500000000000000fb3363b11c",
    x"030b0000000000000155fffffffffffff50003ea0f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2d01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f338f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13b41c",
    x"070a0000000000000155fffffffffffff8ef35ef9f1c",
    x"08020000000000000155fffffffffffff6f669dcc31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec921c",
    x"0209000000000000015500000000000000fb3363ab1c",
    x"030b0000000000000155fffffffffffff50003ea101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2cd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f338b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13ad1c",
    x"070a0000000000000155fffffffffffff8ef35ef9c1c",
    x"08020000000000000155fffffffffffff6f669dcc11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec931c",
    x"0209000000000000015500000000000000fb3363a61c",
    x"030b0000000000000155fffffffffffff50003ea111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2cb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13a71c",
    x"070a0000000000000155fffffffffffff8ef35ef981c",
    x"08020000000000000155fffffffffffff6f669dcbf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec941c",
    x"0209000000000000015500000000000000fb3363a01c",
    x"030b0000000000000155fffffffffffff50003ea121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2c81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13a11c",
    x"070a0000000000000155fffffffffffff8ef35ef941c",
    x"08020000000000000155fffffffffffff6f669dcbc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec951c",
    x"0209000000000000015500000000000000fb33639b1c",
    x"030b0000000000000155fffffffffffff50003ea121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2c61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd139b1c",
    x"070a0000000000000155fffffffffffff8ef35ef901c",
    x"08020000000000000155fffffffffffff6f669dcba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec961c",
    x"0209000000000000015500000000000000fb3363951c",
    x"030b0000000000000155fffffffffffff50003ea131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2c31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f337d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13951c",
    x"070a0000000000000155fffffffffffff8ef35ef8d1c",
    x"08020000000000000155fffffffffffff6f669dcb71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec971c",
    x"0209000000000000015500000000000000fb33638f1c",
    x"030b0000000000000155fffffffffffff50003ea141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2c11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd138f1c",
    x"070a0000000000000155fffffffffffff8ef35ef891c",
    x"08020000000000000155fffffffffffff6f669dcb51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec981c",
    x"0209000000000000015500000000000000fb33638a1c",
    x"030b0000000000000155fffffffffffff50003ea151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2be1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13881c",
    x"070a0000000000000155fffffffffffff8ef35ef851c",
    x"08020000000000000155fffffffffffff6f669dcb31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c7b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbec991c",
    x"0209000000000000025500000000000000fb3363841c",
    x"030b0000000000000255fffffffffffff50003ea161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dc2bc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f33721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd13821c",
    x"070a0000000000000255fffffffffffff8ef35ef821c",
    x"08020000000000000255fffffffffffff6f669dcb01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbec9b1c",
    x"0209000000000000015500000000000000fb33637e1c",
    x"030b0000000000000155fffffffffffff50003ea171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2b91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f336e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd137c1c",
    x"070a0000000000000155fffffffffffff8ef35ef7e1c",
    x"08020000000000000155fffffffffffff6f669dcae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c7aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbec9c1c",
    x"0209000000000000031f00000000000000fb3363791c",
    x"030b000000000000031ffffffffffffff50003ea181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc2b71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f336b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd13761c",
    x"070a000000000000031ffffffffffffff8ef35ef7a1c",
    x"0802000000000000031ffffffffffffff6f669dcab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c7a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbec9d1c",
    x"020900000000000000ae00000000000000fb3363731c",
    x"030b00000000000000aefffffffffffff50003ea191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc2b41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f33671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd13701c",
    x"070a00000000000000aefffffffffffff8ef35ef761c",
    x"080200000000000000aefffffffffffff6f669dca91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c7a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbec9e1c",
    x"020900000000000001a400000000000000fb33636e1c",
    x"030b00000000000001a4fffffffffffff50003ea1a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc2b21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f33641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd13691c",
    x"070a00000000000001a4fffffffffffff8ef35ef731c",
    x"080200000000000001a4fffffffffffff6f669dca61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266c79d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbec9f1c",
    x"0209000000000000019600000000000000fb3363681c",
    x"030b0000000000000196fffffffffffff50003ea1a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc2af1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f33601c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001960000000000000004cd13631c",
    x"070a0000000000000196fffffffffffff8ef35ef6f1c",
    x"08020000000000000196fffffffffffff6f669dca41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca01c",
    x"0209000000000000015500000000000000fb3363621c",
    x"030b0000000000000155fffffffffffff50003ea1b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2ad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f335c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd135d1c",
    x"070a0000000000000155fffffffffffff8ef35ef6b1c",
    x"08020000000000000155fffffffffffff6f669dca21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca11c",
    x"0209000000000000015500000000000000fb33635d1c",
    x"030b0000000000000155fffffffffffff50003ea1c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2aa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13571c",
    x"070a0000000000000155fffffffffffff8ef35ef671c",
    x"08020000000000000155fffffffffffff6f669dc9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca31c",
    x"0209000000000000015500000000000000fb3363571c",
    x"030b0000000000000155fffffffffffff50003ea1d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2a81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13511c",
    x"070a0000000000000155fffffffffffff8ef35ef641c",
    x"08020000000000000155fffffffffffff6f669dc9d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c78c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca41c",
    x"0209000000000000015500000000000000fb3363521c",
    x"030b0000000000000155fffffffffffff50003ea1e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2a51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd134b1c",
    x"070a0000000000000155fffffffffffff8ef35ef601c",
    x"08020000000000000155fffffffffffff6f669dc9a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca51c",
    x"0209000000000000015500000000000000fb33634c1c",
    x"030b0000000000000155fffffffffffff50003ea1f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2a31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f334e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13441c",
    x"070a0000000000000155fffffffffffff8ef35ef5c1c",
    x"08020000000000000155fffffffffffff6f669dc981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca61c",
    x"0209000000000000015500000000000000fb3363461c",
    x"030b0000000000000155fffffffffffff50003ea201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2a01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f334a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd133e1c",
    x"070a0000000000000155fffffffffffff8ef35ef591c",
    x"08020000000000000155fffffffffffff6f669dc961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca71c",
    x"0209000000000000015500000000000000fb3363411c",
    x"030b0000000000000155fffffffffffff50003ea211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc29e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13381c",
    x"070a0000000000000155fffffffffffff8ef35ef551c",
    x"08020000000000000155fffffffffffff6f669dc931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c77c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca81c",
    x"0209000000000000015500000000000000fb33633b1c",
    x"030b0000000000000155fffffffffffff50003ea221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc29b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33431c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13321c",
    x"070a0000000000000155fffffffffffff8ef35ef511c",
    x"08020000000000000155fffffffffffff6f669dc911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeca91c",
    x"0209000000000000015500000000000000fb3363351c",
    x"030b0000000000000155fffffffffffff50003ea221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2981c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd132c1c",
    x"070a0000000000000155fffffffffffff8ef35ef4d1c",
    x"08020000000000000155fffffffffffff6f669dc8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecab1c",
    x"0209000000000000015500000000000000fb3363301c",
    x"030b0000000000000155fffffffffffff50003ea231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2961c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f333c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13251c",
    x"070a0000000000000155fffffffffffff8ef35ef4a1c",
    x"08020000000000000155fffffffffffff6f669dc8c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c76f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecac1c",
    x"0209000000000000015500000000000000fb33632a1c",
    x"030b0000000000000155fffffffffffff50003ea241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2931c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33381c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd131f1c",
    x"070a0000000000000155fffffffffffff8ef35ef461c",
    x"08020000000000000155fffffffffffff6f669dc891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c76b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecad1c",
    x"0209000000000000015500000000000000fb3363251c",
    x"030b0000000000000155fffffffffffff50003ea251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13191c",
    x"070a0000000000000155fffffffffffff8ef35ef421c",
    x"08020000000000000155fffffffffffff6f669dc871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecae1c",
    x"0209000000000000015500000000000000fb33631f1c",
    x"030b0000000000000155fffffffffffff50003ea261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc28e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33311c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd13131c",
    x"070a0000000000000155fffffffffffff8ef35ef3f1c",
    x"08020000000000000155fffffffffffff6f669dc851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecaf1c",
    x"0209000000000000015500000000000000fb3363191c",
    x"030b0000000000000155fffffffffffff50003ea271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc28c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f332d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd130d1c",
    x"070a0000000000000155fffffffffffff8ef35ef3b1c",
    x"08020000000000000155fffffffffffff6f669dc821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266c75f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbecb01c",
    x"020900000000000002a500000000000000fb3363141c",
    x"030b00000000000002a5fffffffffffff50003ea281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc2891c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f332a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd13071c",
    x"070a00000000000002a5fffffffffffff8ef35ef371c",
    x"080200000000000002a5fffffffffffff6f669dc801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c75a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecb11c",
    x"020900000000000002aa00000000000000fb33630e1c",
    x"030b00000000000002aafffffffffffff50003ea291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33261c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd13001c",
    x"070a00000000000002aafffffffffffff8ef35ef331c",
    x"080200000000000002aafffffffffffff6f669dc7d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c7561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbecb21c",
    x"0209000000000000031f00000000000000fb3363081c",
    x"030b000000000000031ffffffffffffff50003ea2a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc2841c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f33231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd12fa1c",
    x"070a000000000000031ffffffffffffff8ef35ef301c",
    x"0802000000000000031ffffffffffffff6f669dc7b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c7521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbecb41c",
    x"020900000000000000ae00000000000000fb3363031c",
    x"030b00000000000000aefffffffffffff50003ea2a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc2821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f331f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd12f41c",
    x"070a00000000000000aefffffffffffff8ef35ef2c1c",
    x"080200000000000000aefffffffffffff6f669dc791c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c74e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbecb51c",
    x"020900000000000001a400000000000000fb3362fd1c",
    x"030b00000000000001a4fffffffffffff50003ea2b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc27f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f331b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd12ee1c",
    x"070a00000000000001a4fffffffffffff8ef35ef281c",
    x"080200000000000001a4fffffffffffff6f669dc761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266c74a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbecb61c",
    x"020900000000000002a600000000000000fb3362f81c",
    x"030b00000000000002a6fffffffffffff50003ea2c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc27d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f33181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd12e81c",
    x"070a00000000000002a6fffffffffffff8ef35ef241c",
    x"080200000000000002a6fffffffffffff6f669dc741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c7461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecb71c",
    x"020900000000000002aa00000000000000fb3362f21c",
    x"030b00000000000002aafffffffffffff50003ea2d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc27a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f33141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd12e11c",
    x"070a00000000000002aafffffffffffff8ef35ef211c",
    x"080200000000000002aafffffffffffff6f669dc711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266c7421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbecb81c",
    x"0209000000000000016900000000000000fb3362ec1c",
    x"030b0000000000000169fffffffffffff50003ea2e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dc2781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001690000000000000b072f33111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd12db1c",
    x"070a0000000000000169fffffffffffff8ef35ef1d1c",
    x"08020000000000000169fffffffffffff6f669dc6f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c73d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecb91c",
    x"0209000000000000015500000000000000fb3362e71c",
    x"030b0000000000000155fffffffffffff50003ea2f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f330d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12d51c",
    x"070a0000000000000155fffffffffffff8ef35ef191c",
    x"08020000000000000155fffffffffffff6f669dc6c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecba1c",
    x"0209000000000000015500000000000000fb3362e11c",
    x"030b0000000000000155fffffffffffff50003ea301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12cf1c",
    x"070a0000000000000155fffffffffffff8ef35ef161c",
    x"08020000000000000155fffffffffffff6f669dc6a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecbc1c",
    x"0209000000000000015500000000000000fb3362dc1c",
    x"030b0000000000000155fffffffffffff50003ea311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12c91c",
    x"070a0000000000000155fffffffffffff8ef35ef121c",
    x"08020000000000000155fffffffffffff6f669dc681c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecbd1c",
    x"0209000000000000015500000000000000fb3362d61c",
    x"030b0000000000000155fffffffffffff50003ea321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc26e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f33021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12c21c",
    x"070a0000000000000155fffffffffffff8ef35ef0e1c",
    x"08020000000000000155fffffffffffff6f669dc651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c72d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecbe1c",
    x"0209000000000000015500000000000000fb3362d01c",
    x"030b0000000000000155fffffffffffff50003ea321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc26b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12bc1c",
    x"070a0000000000000155fffffffffffff8ef35ef0a1c",
    x"08020000000000000155fffffffffffff6f669dc631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7291c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecbf1c",
    x"0209000000000000015500000000000000fb3362cb1c",
    x"030b0000000000000155fffffffffffff50003ea331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32fb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12b61c",
    x"070a0000000000000155fffffffffffff8ef35ef071c",
    x"08020000000000000155fffffffffffff6f669dc601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecc01c",
    x"0209000000000000015500000000000000fb3362c51c",
    x"030b0000000000000155fffffffffffff50003ea341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32f71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12b01c",
    x"070a0000000000000155fffffffffffff8ef35ef031c",
    x"08020000000000000155fffffffffffff6f669dc5e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecc11c",
    x"0209000000000000015500000000000000fb3362bf1c",
    x"030b0000000000000155fffffffffffff50003ea351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12aa1c",
    x"070a0000000000000155fffffffffffff8ef35eeff1c",
    x"08020000000000000155fffffffffffff6f669dc5b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c71c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecc21c",
    x"0209000000000000015500000000000000fb3362ba1c",
    x"030b0000000000000155fffffffffffff50003ea361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32f01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12a41c",
    x"070a0000000000000155fffffffffffff8ef35eefc1c",
    x"08020000000000000155fffffffffffff6f669dc591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecc41c",
    x"0209000000000000015500000000000000fb3362b41c",
    x"030b0000000000000155fffffffffffff50003ea371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc25f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd129d1c",
    x"070a0000000000000155fffffffffffff8ef35eef81c",
    x"08020000000000000155fffffffffffff6f669dc571c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecc51c",
    x"0209000000000000015500000000000000fb3362af1c",
    x"030b0000000000000155fffffffffffff50003ea381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc25c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32e91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12971c",
    x"070a0000000000000155fffffffffffff8ef35eef41c",
    x"08020000000000000155fffffffffffff6f669dc541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c7101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecc61c",
    x"0209000000000000015500000000000000fb3362a91c",
    x"030b0000000000000155fffffffffffff50003ea391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc25a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32e51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12911c",
    x"070a0000000000000155fffffffffffff8ef35eef01c",
    x"08020000000000000155fffffffffffff6f669dc521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266c70b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbecc71c",
    x"0209000000000000019500000000000000fb3362a31c",
    x"030b0000000000000195fffffffffffff50003ea3a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dc2571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f32e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001950000000000000004cd128b1c",
    x"070a0000000000000195fffffffffffff8ef35eeed1c",
    x"08020000000000000195fffffffffffff6f669dc4f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c7071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecc81c",
    x"020900000000000002aa00000000000000fb33629e1c",
    x"030b00000000000002aafffffffffffff50003ea3a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32de1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd12851c",
    x"070a00000000000002aafffffffffffff8ef35eee91c",
    x"080200000000000002aafffffffffffff6f669dc4d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c7031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbecc91c",
    x"0209000000000000031f00000000000000fb3362981c",
    x"030b000000000000031ffffffffffffff50003ea3b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc2521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f32db1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd127e1c",
    x"070a000000000000031ffffffffffffff8ef35eee51c",
    x"0802000000000000031ffffffffffffff6f669dc4b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c6ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbecca1c",
    x"020900000000000000ae00000000000000fb3362931c",
    x"030b00000000000000aefffffffffffff50003ea3c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc24f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f32d71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd12781c",
    x"070a00000000000000aefffffffffffff8ef35eee11c",
    x"080200000000000000aefffffffffffff6f669dc481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c6fb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbeccc1c",
    x"020900000000000001a400000000000000fb33628d1c",
    x"030b00000000000001a4fffffffffffff50003ea3d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc24d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f32d31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd12721c",
    x"070a00000000000001a4fffffffffffff8ef35eede1c",
    x"080200000000000001a4fffffffffffff6f669dc461c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266c6f71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbeccd1c",
    x"020900000000000001a600000000000000fb3362871c",
    x"030b00000000000001a6fffffffffffff50003ea3e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc24a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f32d01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd126c1c",
    x"070a00000000000001a6fffffffffffff8ef35eeda1c",
    x"080200000000000001a6fffffffffffff6f669dc431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6f21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecce1c",
    x"0209000000000000015500000000000000fb3362821c",
    x"030b0000000000000155fffffffffffff50003ea3f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2481c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32cc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12661c",
    x"070a0000000000000155fffffffffffff8ef35eed61c",
    x"08020000000000000155fffffffffffff6f669dc411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeccf1c",
    x"0209000000000000015500000000000000fb33627c1c",
    x"030b0000000000000155fffffffffffff50003ea401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12601c",
    x"070a0000000000000155fffffffffffff8ef35eed31c",
    x"08020000000000000155fffffffffffff6f669dc3e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6ea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd01c",
    x"0209000000000000015500000000000000fb3362761c",
    x"030b0000000000000155fffffffffffff50003ea411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2431c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32c51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12591c",
    x"070a0000000000000155fffffffffffff8ef35eecf1c",
    x"08020000000000000155fffffffffffff6f669dc3c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6e61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd11c",
    x"0209000000000000015500000000000000fb3362711c",
    x"030b0000000000000155fffffffffffff50003ea421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2401c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32c11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12531c",
    x"070a0000000000000155fffffffffffff8ef35eecb1c",
    x"08020000000000000155fffffffffffff6f669dc3a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6e21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd21c",
    x"0209000000000000015500000000000000fb33626b1c",
    x"030b0000000000000155fffffffffffff50003ea421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc23e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd124d1c",
    x"070a0000000000000155fffffffffffff8ef35eec71c",
    x"08020000000000000155fffffffffffff6f669dc371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6de1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd31c",
    x"0209000000000000015500000000000000fb3362661c",
    x"030b0000000000000155fffffffffffff50003ea431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc23b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32ba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12471c",
    x"070a0000000000000155fffffffffffff9ef35eec41c",
    x"08020000000000000155fffffffffffff6f669dc351c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6da1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd51c",
    x"0209000000000000015500000000000000fb3362601c",
    x"030b0000000000000155fffffffffffff50003ea441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12411c",
    x"070a0000000000000155fffffffffffff9ef35eec01c",
    x"08020000000000000155fffffffffffff6f669dc321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6d51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd61c",
    x"0209000000000000015500000000000000fb33625a1c",
    x"030b0000000000000155fffffffffffff50003ea451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32b31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd123a1c",
    x"070a0000000000000155fffffffffffff9ef35eebc1c",
    x"08020000000000000155fffffffffffff6f669dc301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6d11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd71c",
    x"0209000000000000015500000000000000fb3362551c",
    x"030b0000000000000155fffffffffffff50003ea461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32af1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12341c",
    x"070a0000000000000155fffffffffffff9ef35eeb91c",
    x"08020000000000000155fffffffffffff6f669dc2e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6cd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd81c",
    x"0209000000000000015500000000000000fb33624f1c",
    x"030b0000000000000155fffffffffffff50003ea471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd122e1c",
    x"070a0000000000000155fffffffffffff9ef35eeb51c",
    x"08020000000000000155fffffffffffff6f669dc2b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6c91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecd91c",
    x"0209000000000000015500000000000000fb3362491c",
    x"030b0000000000000155fffffffffffff50003ea481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc22f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32a81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12281c",
    x"070a0000000000000155fffffffffffff9ef35eeb11c",
    x"08020000000000000155fffffffffffff6f669dc291c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6c51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecda1c",
    x"0209000000000000015500000000000000fb3362441c",
    x"030b0000000000000155fffffffffffff50003ea491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc22c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12221c",
    x"070a0000000000000155fffffffffffff9ef35eead1c",
    x"08020000000000000155fffffffffffff6f669dc261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6c11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecdb1c",
    x"0209000000000000015500000000000000fb33623e1c",
    x"030b0000000000000155fffffffffffff50003ea4a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc22a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32a11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd121c1c",
    x"070a0000000000000155fffffffffffff9ef35eeaa1c",
    x"08020000000000000155fffffffffffff6f669dc241c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6bc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecdd1c",
    x"0209000000000000015500000000000000fb3362391c",
    x"030b0000000000000155fffffffffffff50003ea4a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2271c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f329d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd12151c",
    x"070a0000000000000155fffffffffffff9ef35eea61c",
    x"08020000000000000155fffffffffffff6f669dc211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c6b81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbecde1c",
    x"0209000000000000029500000000000000fb3362331c",
    x"030b0000000000000295fffffffffffff50003ea4b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc2251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f329a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd120f1c",
    x"070a0000000000000295fffffffffffff9ef35eea21c",
    x"08020000000000000295fffffffffffff6f669dc1f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6b41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecdf1c",
    x"020900000000000002aa00000000000000fb33622d1c",
    x"030b00000000000002aafffffffffffff50003ea4c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc2221c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd12091c",
    x"070a00000000000002aafffffffffffff9ef35ee9e1c",
    x"080200000000000002aafffffffffffff6f669dc1d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c6b01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbece01c",
    x"0209000000000000031f00000000000000fb3362281c",
    x"030b000000000000031ffffffffffffff50003ea4d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc2201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f32931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd12031c",
    x"070a000000000000031ffffffffffffff9ef35ee9b1c",
    x"0802000000000000031ffffffffffffff6f669dc1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c6ac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbece11c",
    x"020900000000000000ae00000000000000fb3362221c",
    x"030b00000000000000aefffffffffffff50003ea4e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc21d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f328f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd11fd1c",
    x"070a00000000000000aefffffffffffff9ef35ee971c",
    x"080200000000000000aefffffffffffff6f669dc181c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c6a81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbece21c",
    x"020900000000000001a400000000000000fb33621d1c",
    x"030b00000000000001a4fffffffffffff50003ea4f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc21b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f328b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd11f61c",
    x"070a00000000000001a4fffffffffffff9ef35ee931c",
    x"080200000000000001a4fffffffffffff6f669dc151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266c6a31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbece31c",
    x"0209000000000000016600000000000000fb3362171c",
    x"030b0000000000000166fffffffffffff50003ea501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc2181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f32881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd11f01c",
    x"070a0000000000000166fffffffffffff9ef35ee901c",
    x"08020000000000000166fffffffffffff6f669dc131c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c69f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbece51c",
    x"0209000000000000015500000000000000fb3362111c",
    x"030b0000000000000155fffffffffffff50003ea511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2151c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11ea1c",
    x"070a0000000000000155fffffffffffff9ef35ee8c1c",
    x"08020000000000000155fffffffffffff6f669dc101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000165ffffffffffffff0266c69b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbece61c",
    x"0209000000000000016500000000000000fb33620c1c",
    x"030b0000000000000165fffffffffffff50003ea511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc2131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f32811c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd11e41c",
    x"070a0000000000000165fffffffffffff9ef35ee881c",
    x"08020000000000000165fffffffffffff6f669dc0e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6971c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbece71c",
    x"0209000000000000015500000000000000fb3362061c",
    x"030b0000000000000155fffffffffffff50003ea521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2101c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f327d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11de1c",
    x"070a0000000000000155fffffffffffff9ef35ee841c",
    x"08020000000000000155fffffffffffff6f669dc0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbece81c",
    x"0209000000000000015500000000000000fb3362001c",
    x"030b0000000000000155fffffffffffff50003ea531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc20e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11d71c",
    x"070a0000000000000155fffffffffffff9ef35ee811c",
    x"08020000000000000155fffffffffffff6f669dc091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c68f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbece91c",
    x"0209000000000000015500000000000000fb3361fb1c",
    x"030b0000000000000155fffffffffffff50003ea541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc20b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11d11c",
    x"070a0000000000000155fffffffffffff9ef35ee7d1c",
    x"08020000000000000155fffffffffffff6f669dc071c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c68a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecea1c",
    x"0209000000000000015500000000000000fb3361f51c",
    x"030b0000000000000155fffffffffffff50003ea551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11cb1c",
    x"070a0000000000000155fffffffffffff9ef35ee791c",
    x"08020000000000000155fffffffffffff6f669dc041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6861c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeceb1c",
    x"0209000000000000015500000000000000fb3361f01c",
    x"030b0000000000000155fffffffffffff50003ea561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2061c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f326f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11c51c",
    x"070a0000000000000155fffffffffffff9ef35ee751c",
    x"08020000000000000155fffffffffffff6f669dc021c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6821c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeced1c",
    x"0209000000000000015500000000000000fb3361ea1c",
    x"030b0000000000000155fffffffffffff50003ea571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f326b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11bf1c",
    x"070a0000000000000155fffffffffffff9ef35ee721c",
    x"08020000000000000155fffffffffffff6f669dc001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c67e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecee1c",
    x"0209000000000000015500000000000000fb3361e41c",
    x"030b0000000000000155fffffffffffff50003ea581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc2011c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11b91c",
    x"070a0000000000000155fffffffffffff9ef35ee6e1c",
    x"08020000000000000155fffffffffffff6f669dbfd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c67a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecef1c",
    x"0209000000000000015500000000000000fb3361df1c",
    x"030b0000000000000155fffffffffffff50003ea591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1ff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11b21c",
    x"070a0000000000000155fffffffffffff9ef35ee6a1c",
    x"08020000000000000155fffffffffffff6f669dbfb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecf01c",
    x"0209000000000000015500000000000000fb3361d91c",
    x"030b0000000000000155fffffffffffff50003ea591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1fc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32601c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11ac1c",
    x"070a0000000000000155fffffffffffff9ef35ee671c",
    x"08020000000000000155fffffffffffff6f669dbf81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecf11c",
    x"0209000000000000015500000000000000fb3361d31c",
    x"030b0000000000000155fffffffffffff50003ea5a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1fa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f325d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11a61c",
    x"070a0000000000000155fffffffffffff9ef35ee631c",
    x"08020000000000000155fffffffffffff6f669dbf61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c66d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecf21c",
    x"0209000000000000015500000000000000fb3361ce1c",
    x"030b0000000000000155fffffffffffff50003ea5b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1f71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd11a01c",
    x"070a0000000000000155fffffffffffff9ef35ee5f1c",
    x"08020000000000000155fffffffffffff6f669dbf31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c6691c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbecf31c",
    x"0209000000000000015500000000000000fb3361c81c",
    x"030b0000000000000155fffffffffffff50003ea5c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1f51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f32551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd119a1c",
    x"070a0000000000000155fffffffffffff9ef35ee5b1c",
    x"08020000000000000155fffffffffffff6f669dbf11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c6651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbecf51c",
    x"0209000000000000025500000000000000fb3361c31c",
    x"030b0000000000000255fffffffffffff50003ea5d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dc1f21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f32521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd11931c",
    x"070a0000000000000255fffffffffffff9ef35ee581c",
    x"08020000000000000255fffffffffffff6f669dbef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecf61c",
    x"020900000000000002aa00000000000000fb3361bd1c",
    x"030b00000000000002aafffffffffffff50003ea5e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1f01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f324e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd118d1c",
    x"070a00000000000002aafffffffffffff9ef35ee541c",
    x"080200000000000002aafffffffffffff6f669dbec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c65d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbecf71c",
    x"0209000000000000031f00000000000000fb3361b71c",
    x"030b000000000000031ffffffffffffff50003ea5f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc1ed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f324b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd11871c",
    x"070a000000000000031ffffffffffffff9ef35ee501c",
    x"0802000000000000031ffffffffffffff6f669dbea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c6591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbecf81c",
    x"020900000000000000ae00000000000000fb3361b21c",
    x"030b00000000000000aefffffffffffff50003ea601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc1eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f32471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd11811c",
    x"070a00000000000000aefffffffffffff9ef35ee4c1c",
    x"080200000000000000aefffffffffffff6f669dbe71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c6541c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbecf91c",
    x"020900000000000001a400000000000000fb3361ac1c",
    x"030b00000000000001a4fffffffffffff50003ea601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc1e81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f32431c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd117b1c",
    x"070a00000000000001a4fffffffffffff9ef35ee491c",
    x"080200000000000001a4fffffffffffff6f669dbe51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266c6501c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbecfa1c",
    x"0209000000000000026600000000000000fb3361a71c",
    x"030b0000000000000266fffffffffffff50003ea611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc1e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f32401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002660000000000000004cd11751c",
    x"070a0000000000000266fffffffffffff9ef35ee451c",
    x"08020000000000000266fffffffffffff6f669dbe31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c64c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecfb1c",
    x"020900000000000002aa00000000000000fb3361a11c",
    x"030b00000000000002aafffffffffffff50003ea621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1e31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f323c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd116e1c",
    x"070a00000000000002aafffffffffffff9ef35ee411c",
    x"080200000000000002aafffffffffffff6f669dbe01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecfc1c",
    x"020900000000000002aa00000000000000fb33619b1c",
    x"030b00000000000002aafffffffffffff50003ea631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11681c",
    x"070a00000000000002aafffffffffffff9ef35ee3e1c",
    x"080200000000000002aafffffffffffff6f669dbde1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecfe1c",
    x"020900000000000002aa00000000000000fb3361961c",
    x"030b00000000000002aafffffffffffff50003ea641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1de1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11621c",
    x"070a00000000000002aafffffffffffff9ef35ee3a1c",
    x"080200000000000002aafffffffffffff6f669dbdb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbecff1c",
    x"020900000000000002aa00000000000000fb3361901c",
    x"030b00000000000002aafffffffffffff50003ea651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1db1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32311c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd115c1c",
    x"070a00000000000002aafffffffffffff9ef35ee361c",
    x"080200000000000002aafffffffffffff6f669dbd91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c63b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed001c",
    x"020900000000000002aa00000000000000fb33618a1c",
    x"030b00000000000002aafffffffffffff50003ea661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1d91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f322e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11561c",
    x"070a00000000000002aafffffffffffff9ef35ee321c",
    x"080200000000000002aafffffffffffff6f669dbd61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6371c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed011c",
    x"020900000000000002aa00000000000000fb3361851c",
    x"030b00000000000002aafffffffffffff50003ea671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1d61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f322a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd114f1c",
    x"070a00000000000002aafffffffffffff9ef35ee2f1c",
    x"080200000000000002aafffffffffffff6f669dbd41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6331c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed021c",
    x"020900000000000002aa00000000000000fb33617f1c",
    x"030b00000000000002aafffffffffffff50003ea681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1d41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11491c",
    x"070a00000000000002aafffffffffffff9ef35ee2b1c",
    x"080200000000000002aafffffffffffff6f669dbd21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c62f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed031c",
    x"020900000000000002aa00000000000000fb33617a1c",
    x"030b00000000000002aafffffffffffff50003ea681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1d11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11431c",
    x"070a00000000000002aafffffffffffff9ef35ee271c",
    x"080200000000000002aafffffffffffff6f669dbcf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c62b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed041c",
    x"020900000000000002aa00000000000000fb3361741c",
    x"030b00000000000002aafffffffffffff50003ea691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1cf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd113d1c",
    x"070a00000000000002aafffffffffffff9ef35ee231c",
    x"080200000000000002aafffffffffffff6f669dbcd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed061c",
    x"020900000000000002aa00000000000000fb33616e1c",
    x"030b00000000000002aafffffffffffff50003ea6a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1cc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f321c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11371c",
    x"070a00000000000002aafffffffffffff9ef35ee201c",
    x"080200000000000002aafffffffffffff6f669dbca1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed071c",
    x"020900000000000002aa00000000000000fb3361691c",
    x"030b00000000000002aafffffffffffff50003ea6b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1ca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32181c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11301c",
    x"070a00000000000002aafffffffffffff9ef35ee1c1c",
    x"080200000000000002aafffffffffffff6f669dbc81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c61e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed081c",
    x"020900000000000002aa00000000000000fb3361631c",
    x"030b00000000000002aafffffffffffff50003ea6c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1c71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd112a1c",
    x"070a00000000000002aafffffffffffff9ef35ee181c",
    x"080200000000000002aafffffffffffff6f669dbc51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c61a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed091c",
    x"020900000000000002aa00000000000000fb33615d1c",
    x"030b00000000000002aafffffffffffff50003ea6d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11241c",
    x"070a00000000000002aafffffffffffff9ef35ee141c",
    x"080200000000000002aafffffffffffff6f669dbc31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6161c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed0a1c",
    x"020900000000000002aa00000000000000fb3361581c",
    x"030b00000000000002aafffffffffffff50003ea6e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1c21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f320e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd111e1c",
    x"070a00000000000002aafffffffffffff9ef35ee111c",
    x"080200000000000002aafffffffffffff6f669dbc11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c6121c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed0b1c",
    x"020900000000000002aa00000000000000fb3361521c",
    x"030b00000000000002aafffffffffffff50003ea6f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1c01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f320a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11181c",
    x"070a00000000000002aafffffffffffff9ef35ee0d1c",
    x"080200000000000002aafffffffffffff6f669dbbe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c60e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed0c1c",
    x"020900000000000002aa00000000000000fb33614d1c",
    x"030b00000000000002aafffffffffffff50003ea6f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f32061c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd11121c",
    x"070a00000000000002aafffffffffffff9ef35ee091c",
    x"080200000000000002aafffffffffffff6f669dbbc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c60a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed0e1c",
    x"0209000000000000031f00000000000000fb3361471c",
    x"030b000000000000031ffffffffffffff50003ea701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc1bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f32031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd110b1c",
    x"070a000000000000031ffffffffffffff9ef35ee061c",
    x"0802000000000000031ffffffffffffff6f669dbb91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c6051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed0f1c",
    x"020900000000000000ae00000000000000fb3361411c",
    x"030b00000000000000aefffffffffffff50003ea711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc1b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f31ff1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd11051c",
    x"070a00000000000000aefffffffffffff9ef35ee021c",
    x"080200000000000000aefffffffffffff6f669dbb71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c6011c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed101c",
    x"020900000000000001a400000000000000fb33613c1c",
    x"030b00000000000001a4fffffffffffff50003ea721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc1b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f31fc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd10ff1c",
    x"070a00000000000001a4fffffffffffff9ef35edfe1c",
    x"080200000000000001a4fffffffffffff6f669dbb51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266c5fd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbed111c",
    x"020900000000000001aa00000000000000fb3361361c",
    x"030b00000000000001aafffffffffffff50003ea731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc1b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f31f81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd10f91c",
    x"070a00000000000001aafffffffffffff9ef35edfa1c",
    x"080200000000000001aafffffffffffff6f669dbb21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c5f91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbed121c",
    x"0209000000000000029500000000000000fb3361311c",
    x"030b0000000000000295fffffffffffff50003ea741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc1b11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31f41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd10f31c",
    x"070a0000000000000295fffffffffffff9ef35edf71c",
    x"08020000000000000295fffffffffffff6f669dbb01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266c5f51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbed131c",
    x"0209000000000000015a00000000000000fb33612b1c",
    x"030b000000000000015afffffffffffff50003ea751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc1ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f31f11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd10ec1c",
    x"070a000000000000015afffffffffffff9ef35edf31c",
    x"0802000000000000015afffffffffffff6f669dbad1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266c5f11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbed141c",
    x"0209000000000000019500000000000000fb3361251c",
    x"030b0000000000000195fffffffffffff50003ea761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dc1ab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f31ed1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001950000000000000004cd10e61c",
    x"070a0000000000000195fffffffffffff9ef35edef1c",
    x"08020000000000000195fffffffffffff6f669dbab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266c5ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbed161c",
    x"020900000000000002a900000000000000fb3361201c",
    x"030b0000000000000155fffffffffffff50003ea771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc1a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31ea1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd10e01c",
    x"070a0000000000000155fffffffffffff9ef35edeb1c",
    x"080200000000000002a9fffffffffffff6f669dba81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266c5e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed171c",
    x"0209000000000000029a00000000000000fb33611a1c",
    x"030b0000000000000265fffffffffffff50003ea771c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc1a61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f31e61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd10da1c",
    x"070a0000000000000255fffffffffffff9ef35ede81c",
    x"080200000000000002a9fffffffffffff6f669dba61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c5e41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbed181c",
    x"0209000000000000015a00000000000000fb3361141c",
    x"030b0000000000000265fffffffffffff50003ea781c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc1a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f31e21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd10d41c",
    x"070a000000000000029afffffffffffff9ef35ede41c",
    x"0802000000000000019afffffffffffff6f669dba41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a9ffffffffffffff0266c5e01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbed191c",
    x"0209000000000000019900000000000000fb33610f1c",
    x"030b0000000000000166fffffffffffff50003ea791c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc1a11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f31df1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd10cd1c",
    x"070a00000000000001a9fffffffffffff9ef35ede01c",
    x"0802000000000000026afffffffffffff6f669dba11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266c5dc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002690000000000000b0bfbed1a1c",
    x"0209000000000000016600000000000000fb3361091c",
    x"030b00000000000001a6fffffffffffff50003ea7a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc19f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f31db1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd10c71c",
    x"070a0000000000000199fffffffffffff9ef35eddd1c",
    x"0802000000000000025afffffffffffff6f669db9f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266c5d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed1b1c",
    x"0209000000000000015500000000000000fb3361041c",
    x"030b000000000000015afffffffffffff50003ea7b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc19c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f31d81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd10c11c",
    x"070a000000000000016afffffffffffff9ef35edd91c",
    x"0802000000000000025afffffffffffff6f669db9c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266c5d41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbed1c1c",
    x"0209000000000000015a00000000000000fb3360fe1c",
    x"030b0000000000000295fffffffffffff50003ea7c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc19a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f31d41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd10bb1c",
    x"070a00000000000001aafffffffffffff9ef35edd51c",
    x"08020000000000000296fffffffffffff6f669db9a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266c5cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002990000000000000b0bfbed1e1c",
    x"020900000000000001a900000000000000fb3360f81c",
    x"030b0000000000000299fffffffffffff50003ea7d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dc1971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f31d01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd10b51c",
    x"070a0000000000000165fffffffffffff9ef35edd11c",
    x"0802000000000000016afffffffffffff6f669db971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266c5cb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbed1f1c",
    x"020900000000000002aa00000000000000fb3360f31c",
    x"030b0000000000000169fffffffffffff50003ea7e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc1951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31cd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd10af1c",
    x"070a00000000000002a9fffffffffffff9ef35edce1c",
    x"08020000000000000199fffffffffffff6f669db951c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000299ffffffffffffff0266c5c71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbed201c",
    x"0209000000000000029a00000000000000fb3360ed1c",
    x"030b000000000000019afffffffffffff50003ea7e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc1921c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31c91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd10a81c",
    x"070a000000000000016afffffffffffff9ef35edca1c",
    x"08020000000000000165fffffffffffff6f669db931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266c5c31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbed211c",
    x"020900000000000002a600000000000000fb3360e71c",
    x"030b000000000000015afffffffffffff50003ea7f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc1901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31c61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd10a21c",
    x"070a000000000000025afffffffffffff9ef35edc61c",
    x"0802000000000000025afffffffffffff6f669db901c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266c5bf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbed221c",
    x"0209000000000000016a00000000000000fb3360e21c",
    x"030b00000000000001a5fffffffffffff50003ea801c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc18d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f31c21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd109c1c",
    x"070a0000000000000299fffffffffffff9ef35edc21c",
    x"08020000000000000269fffffffffffff6f669db8e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266c5bb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbed231c",
    x"020900000000000002a600000000000000fb3360dc1c",
    x"030b0000000000000159fffffffffffff50003ea811c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc18b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f31be1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd10961c",
    x"070a0000000000000159fffffffffffff9ef35edbf1c",
    x"08020000000000000295fffffffffffff6f669db8b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c5b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed241c",
    x"0209000000000000031f00000000000000fb3360d71c",
    x"030b000000000000031ffffffffffffff50003ea821c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc1881c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f31bb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd10901c",
    x"070a000000000000031ffffffffffffff9ef35edbb1c",
    x"0802000000000000031ffffffffffffff6f669db891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c5b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed261c",
    x"020900000000000000ae00000000000000fb3360d11c",
    x"030b00000000000000aefffffffffffff50003ea831c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc1861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f31b71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd10891c",
    x"070a00000000000000aefffffffffffff9ef35edb71c",
    x"080200000000000000aefffffffffffff6f669db871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c5ae1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed271c",
    x"020900000000000001a400000000000000fb3360cb1c",
    x"030b00000000000001a4fffffffffffff50003ea841c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc1831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f31b41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd10831c",
    x"070a00000000000001a4fffffffffffff9ef35edb31c",
    x"080200000000000001a4fffffffffffff6f669db841c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c5aa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbed281c",
    x"0209000000000000016a00000000000000fb3360c61c",
    x"030b000000000000016afffffffffffff50003ea851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc1801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f31b01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd107d1c",
    x"070a000000000000016afffffffffffff9ef35edb01c",
    x"0802000000000000016afffffffffffff6f669db821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c5a61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed291c",
    x"0209000000000000015500000000000000fb3360c01c",
    x"030b0000000000000155fffffffffffff50003ea851c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc17e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31ac1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd10771c",
    x"070a0000000000000155fffffffffffff9ef35edac1c",
    x"08020000000000000155fffffffffffff6f669db7f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266c5a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbed2a1c",
    x"0209000000000000019500000000000000fb3360bb1c",
    x"030b0000000000000195fffffffffffff50003ea861c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000195fffffffffffff4099dc17b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f31a91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd10711c",
    x"070a0000000000000195fffffffffffff9ef35eda81c",
    x"080200000000000002a5fffffffffffff6f669db7d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c59d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed2b1c",
    x"020900000000000002aa00000000000000fb3360b51c",
    x"030b00000000000002aafffffffffffff50003ea871c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f31a51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd106a1c",
    x"070a00000000000002aafffffffffffff9ef35eda51c",
    x"08020000000000000155fffffffffffff6f669db7a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266c5991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbed2c1c",
    x"0209000000000000029600000000000000fb3360af1c",
    x"030b00000000000001aafffffffffffff50003ea881c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc1761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f31a21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd10641c",
    x"070a0000000000000256fffffffffffff9ef35eda11c",
    x"08020000000000000155fffffffffffff6f669db781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a5ffffffffffffff0266c5951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbed2e1c",
    x"0209000000000000026500000000000000fb3360aa1c",
    x"030b00000000000002a9fffffffffffff50003ea891c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc1741c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f319e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd105e1c",
    x"070a000000000000029afffffffffffff9ef35ed9d1c",
    x"08020000000000000159fffffffffffff6f669db761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266c5911c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbed2f1c",
    x"0209000000000000029600000000000000fb3360a41c",
    x"030b000000000000016afffffffffffff50003ea8a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc1711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f319a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd10581c",
    x"070a0000000000000159fffffffffffff9ef35ed991c",
    x"0802000000000000015afffffffffffff6f669db731c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c58d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed301c",
    x"0209000000000000016900000000000000fb33609e1c",
    x"030b0000000000000295fffffffffffff50003ea8b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc16f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31971c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd10521c",
    x"070a0000000000000196fffffffffffff9ef35ed961c",
    x"08020000000000000299fffffffffffff6f669db711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c5891c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbed311c",
    x"020900000000000002a500000000000000fb3360991c",
    x"030b0000000000000156fffffffffffff50003ea8c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a5fffffffffffff4099dc16c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f31931c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd104c1c",
    x"070a00000000000002a6fffffffffffff9ef35ed921c",
    x"080200000000000001a5fffffffffffff6f669db6e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266c5851c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbed321c",
    x"0209000000000000025500000000000000fb3360931c",
    x"030b000000000000016afffffffffffff50003ea8c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dc16a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f31901c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd10451c",
    x"070a0000000000000295fffffffffffff9ef35ed8e1c",
    x"0802000000000000026afffffffffffff6f669db6c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c5801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbed331c",
    x"0209000000000000029a00000000000000fb33608e1c",
    x"030b0000000000000269fffffffffffff50003ea8d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc1671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f318c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd103f1c",
    x"070a0000000000000196fffffffffffff9ef35ed8a1c",
    x"08020000000000000165fffffffffffff6f669db691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c57c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbed341c",
    x"020900000000000001a600000000000000fb3360881c",
    x"030b000000000000019afffffffffffff50003ea8e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc1651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f31891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd10391c",
    x"070a000000000000026afffffffffffff9ef35ed871c",
    x"0802000000000000019afffffffffffff6f669db671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266c5781c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001990000000000000b0bfbed351c",
    x"0209000000000000025a00000000000000fb3360821c",
    x"030b00000000000002a9fffffffffffff50003ea8f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc1621c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f31851c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a50000000000000004cd10331c",
    x"070a00000000000002a6fffffffffffff9ef35ed831c",
    x"08020000000000000295fffffffffffff6f669db651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266c5741c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbed371c",
    x"0209000000000000029600000000000000fb33607d1c",
    x"030b000000000000025afffffffffffff50003ea901c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000165fffffffffffff4099dc1601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f31811c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd102d1c",
    x"070a000000000000019afffffffffffff9ef35ed7f1c",
    x"0802000000000000029afffffffffffff6f669db621c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266c5701c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbed381c",
    x"0209000000000000019900000000000000fb3360771c",
    x"030b0000000000000156fffffffffffff50003ea911c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dc15d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f317e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd10261c",
    x"070a0000000000000166fffffffffffff9ef35ed7b1c",
    x"080200000000000001a9fffffffffffff6f669db601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c56c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbed391c",
    x"0209000000000000015600000000000000fb3360711c",
    x"030b0000000000000169fffffffffffff50003ea921c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000269fffffffffffff4099dc15b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f317a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd10201c",
    x"070a0000000000000159fffffffffffff9ef35ed781c",
    x"08020000000000000255fffffffffffff6f669db5d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266c5671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed3a1c",
    x"0209000000000000029a00000000000000fb33606c1c",
    x"030b00000000000002a9fffffffffffff50003ea931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc1581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31771c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd101a1c",
    x"070a0000000000000159fffffffffffff9ef35ed741c",
    x"08020000000000000299fffffffffffff6f669db5b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c5631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed3b1c",
    x"0209000000000000031f00000000000000fb3360661c",
    x"030b000000000000031ffffffffffffff50003ea931c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc1561c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f31731c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd10141c",
    x"070a000000000000031ffffffffffffff9ef35ed701c",
    x"0802000000000000031ffffffffffffff6f669db591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c55f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed3c1c",
    x"020900000000000000ae00000000000000fb3360611c",
    x"030b00000000000000aefffffffffffff50003ea941c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc1531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f316f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd100e1c",
    x"070a00000000000000aefffffffffffff9ef35ed6d1c",
    x"080200000000000000aefffffffffffff6f669db561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c55b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed3d1c",
    x"020900000000000001a400000000000000fb33605b1c",
    x"030b00000000000001a4fffffffffffff50003ea951c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc1501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f316c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd10071c",
    x"070a00000000000001a4fffffffffffff9ef35ed691c",
    x"080200000000000001a4fffffffffffff6f669db541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266c5571c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbed3f1c",
    x"0209000000000000026a00000000000000fb3360551c",
    x"030b000000000000026afffffffffffff50003ea961c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc14e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f31681c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026a0000000000000004cd10011c",
    x"070a000000000000026afffffffffffff9ef35ed651c",
    x"0802000000000000026afffffffffffff6f669db511c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c5531c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed401c",
    x"0209000000000000015500000000000000fb3360501c",
    x"030b0000000000000155fffffffffffff50003ea971c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc14b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f31651c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd0ffb1c",
    x"070a00000000000002a9fffffffffffff9ef35ed611c",
    x"08020000000000000155fffffffffffff6f669db4f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c54e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed411c",
    x"0209000000000000015500000000000000fb33604a1c",
    x"030b0000000000000155fffffffffffff50003ea981c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f31611c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ff51c",
    x"070a00000000000001aafffffffffffff9ef35ed5e1c",
    x"08020000000000000155fffffffffffff6f669db4c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266c54a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbed421c",
    x"0209000000000000015600000000000000fb3360441c",
    x"030b0000000000000155fffffffffffff50003ea991c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc1461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f315d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd0fef1c",
    x"070a00000000000002aafffffffffffff9ef35ed5a1c",
    x"08020000000000000155fffffffffffff6f669db4a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c5461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbed431c",
    x"0209000000000000025500000000000000fb33603f1c",
    x"030b0000000000000195fffffffffffff50003ea9a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002690000000000000b072f315a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd0fe91c",
    x"070a000000000000026afffffffffffff9ef35ed561c",
    x"08020000000000000195fffffffffffff6f669db481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266c5421c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbed441c",
    x"0209000000000000016500000000000000fb3360391c",
    x"030b00000000000002a9fffffffffffff50003ea9a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dc1411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31561c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002590000000000000004cd0fe21c",
    x"070a0000000000000256fffffffffffff9ef35ed521c",
    x"08020000000000000299fffffffffffff6f669db451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266c53e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbed451c",
    x"0209000000000000019900000000000000fb3360341c",
    x"030b0000000000000195fffffffffffff50003ea9b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc13f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31531c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd0fdc1c",
    x"070a0000000000000266fffffffffffff9ef35ed4f1c",
    x"080200000000000002a6fffffffffffff6f669db431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266c53a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbed471c",
    x"0209000000000000016500000000000000fb33602e1c",
    x"030b0000000000000166fffffffffffff50003ea9c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dc13c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f314f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd0fd61c",
    x"070a0000000000000156fffffffffffff9ef35ed4b1c",
    x"0802000000000000025afffffffffffff6f669db401c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266c5361c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbed481c",
    x"0209000000000000019500000000000000fb3360281c",
    x"030b0000000000000265fffffffffffff50003ea9d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000199fffffffffffff4099dc13a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f314b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a90000000000000004cd0fd01c",
    x"070a000000000000025afffffffffffff9ef35ed471c",
    x"0802000000000000016afffffffffffff6f669db3e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c5311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbed491c",
    x"0209000000000000026a00000000000000fb3360231c",
    x"030b00000000000002aafffffffffffff50003ea9e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f31481c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd0fca1c",
    x"070a0000000000000195fffffffffffff9ef35ed431c",
    x"08020000000000000195fffffffffffff6f669db3b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000265ffffffffffffff0266c52d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbed4a1c",
    x"0209000000000000025600000000000000fb33601d1c",
    x"030b00000000000002a5fffffffffffff50003ea9f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dc1351c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f31441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd0fc31c",
    x"070a00000000000002a5fffffffffffff9ef35ed401c",
    x"08020000000000000295fffffffffffff6f669db391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c5291c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbed4b1c",
    x"020900000000000001a900000000000000fb3360181c",
    x"030b0000000000000155fffffffffffff50003eaa01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc1321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001650000000000000b072f31411c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd0fbd1c",
    x"070a0000000000000256fffffffffffff9ef35ed3c1c",
    x"08020000000000000199fffffffffffff6f669db371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c5251c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbed4c1c",
    x"0209000000000000029500000000000000fb3360121c",
    x"030b0000000000000299fffffffffffff50003eaa11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1301c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f313d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd0fb71c",
    x"070a0000000000000266fffffffffffff9ef35ed381c",
    x"08020000000000000166fffffffffffff6f669db341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266c5211c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbed4d1c",
    x"0209000000000000016900000000000000fb33600c1c",
    x"030b000000000000016afffffffffffff50003eaa11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc12d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a50000000000000b072f31391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd0fb11c",
    x"070a0000000000000256fffffffffffff9ef35ed341c",
    x"08020000000000000199fffffffffffff6f669db321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266c51d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbed4f1c",
    x"0209000000000000026a00000000000000fb3360071c",
    x"030b000000000000016afffffffffffff50003eaa21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc12a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f31361c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd0fab1c",
    x"070a00000000000001a5fffffffffffff9ef35ed311c",
    x"08020000000000000266fffffffffffff6f669db2f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c5181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbed501c",
    x"020900000000000001a900000000000000fb3360011c",
    x"030b000000000000026afffffffffffff50003eaa31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dc1281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f31321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd0fa41c",
    x"070a0000000000000166fffffffffffff9ef35ed2d1c",
    x"08020000000000000296fffffffffffff6f669db2d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266c5141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbed511c",
    x"020900000000000002a600000000000000fb335ffb1c",
    x"030b000000000000015afffffffffffff50003eaa41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc1251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f312f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002990000000000000004cd0f9e1c",
    x"070a0000000000000295fffffffffffff9ef35ed291c",
    x"080200000000000002a5fffffffffffff6f669db2a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c5101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed521c",
    x"0209000000000000031f00000000000000fb335ff61c",
    x"030b000000000000031ffffffffffffff50003eaa51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc1231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f312b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0f981c",
    x"070a000000000000031ffffffffffffff9ef35ed261c",
    x"0802000000000000031ffffffffffffff6f669db281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c50c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed531c",
    x"020900000000000000ae00000000000000fb335ff01c",
    x"030b00000000000000aefffffffffffff50003eaa61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc1201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f31281c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0f921c",
    x"070a00000000000000aefffffffffffff9ef35ed221c",
    x"080200000000000000aefffffffffffff6f669db261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c5081c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed541c",
    x"020900000000000001a400000000000000fb335feb1c",
    x"030b00000000000001a4fffffffffffff50003eaa71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc11e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f31241c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0f8c1c",
    x"070a00000000000001a4fffffffffffff9ef35ed1e1c",
    x"080200000000000001a4fffffffffffff6f669db231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266c5041c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbed551c",
    x"0209000000000000015a00000000000000fb335fe51c",
    x"030b000000000000015afffffffffffff50003eaa81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dc11b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f31201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd0f861c",
    x"070a000000000000015afffffffffffff9ef35ed1a1c",
    x"0802000000000000015afffffffffffff6f669db211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed571c",
    x"020900000000000001aa00000000000000fb335fdf1c",
    x"030b0000000000000255fffffffffffff50003eaa81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc1191c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f311d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0f7f1c",
    x"070a0000000000000155fffffffffffff9ef35ed171c",
    x"08020000000000000155fffffffffffff6f669db1e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000195ffffffffffffff0266c4fb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001950000000000000b0bfbed581c",
    x"0209000000000000016900000000000000fb335fda1c",
    x"030b0000000000000269fffffffffffff50003eaa91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dc1161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f31191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd0f791c",
    x"070a00000000000002a6fffffffffffff9ef35ed131c",
    x"080200000000000001a5fffffffffffff6f669db1c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000199ffffffffffffff0266c4f71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002650000000000000b0bfbed591c",
    x"020900000000000001a600000000000000fb335fd41c",
    x"030b0000000000000296fffffffffffff50003eaaa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000299fffffffffffff4099dc1141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f31161c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd0f731c",
    x"070a000000000000029afffffffffffff9ef35ed0f1c",
    x"08020000000000000196fffffffffffff6f669db1a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c4f31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbed5a1c",
    x"0209000000000000026900000000000000fb335fce1c",
    x"030b0000000000000255fffffffffffff50003eaab1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc1111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f31121c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001990000000000000004cd0f6d1c",
    x"070a0000000000000265fffffffffffff9ef35ed0b1c",
    x"08020000000000000256fffffffffffff6f669db171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4ef1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbed5b1c",
    x"0209000000000000015600000000000000fb335fc91c",
    x"030b0000000000000155fffffffffffff50003eaac1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc10f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f310e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd0f671c",
    x"070a00000000000002aafffffffffffff9ef35ed081c",
    x"08020000000000000155fffffffffffff6f669db151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c4eb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbed5c1c",
    x"0209000000000000016500000000000000fb335fc31c",
    x"030b0000000000000165fffffffffffff50003eaad1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc10c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f310b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001650000000000000004cd0f601c",
    x"070a000000000000029afffffffffffff9ef35ed041c",
    x"08020000000000000165fffffffffffff6f669db121c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4e71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed5d1c",
    x"020900000000000002aa00000000000000fb335fbe1c",
    x"030b00000000000002aafffffffffffff50003eaae1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc10a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0f5a1c",
    x"070a0000000000000155fffffffffffff9ef35ed001c",
    x"080200000000000002aafffffffffffff6f669db101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4e21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed5f1c",
    x"020900000000000002aa00000000000000fb335fb81c",
    x"030b00000000000002aafffffffffffff50003eaaf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31041c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0f541c",
    x"070a0000000000000155fffffffffffff9ef35ecfc1c",
    x"080200000000000002aafffffffffffff6f669db0d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4de1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed601c",
    x"020900000000000002aa00000000000000fb335fb21c",
    x"030b00000000000002aafffffffffffff50003eaaf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc1041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f31001c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0f4e1c",
    x"070a0000000000000155fffffffffffff9ef35ecf91c",
    x"080200000000000002aafffffffffffff6f669db0b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000259ffffffffffffff0266c4da1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002590000000000000b0bfbed611c",
    x"020900000000000001a600000000000000fb335fad1c",
    x"030b00000000000001a6fffffffffffff50003eab01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000259fffffffffffff4099dc1021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002590000000000000b072f30fc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd0f481c",
    x"070a0000000000000259fffffffffffff9ef35ecf51c",
    x"080200000000000001a6fffffffffffff6f669db091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4d61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed621c",
    x"020900000000000002aa00000000000000fb335fa71c",
    x"030b00000000000002aafffffffffffff50003eab11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0ff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30f91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0f411c",
    x"070a0000000000000155fffffffffffff9ef35ecf11c",
    x"080200000000000002aafffffffffffff6f669db061c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4d21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed631c",
    x"020900000000000002aa00000000000000fb335fa21c",
    x"030b00000000000002aafffffffffffff50003eab21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0fd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30f51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0f3b1c",
    x"070a0000000000000155fffffffffffff9ef35eced1c",
    x"080200000000000002aafffffffffffff6f669db041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c4ce1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbed641c",
    x"020900000000000002a600000000000000fb335f9c1c",
    x"030b00000000000002a6fffffffffffff50003eab31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc0fa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f30f21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd0f351c",
    x"070a0000000000000159fffffffffffff9ef35ecea1c",
    x"080200000000000002a6fffffffffffff6f669db011c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c4c91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a50000000000000b0bfbed651c",
    x"0209000000000000029500000000000000fb335f961c",
    x"030b00000000000002aafffffffffffff50003eab41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dc0f81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001950000000000000b072f30ee1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd0f2f1c",
    x"070a000000000000019afffffffffffff9ef35ece61c",
    x"080200000000000002a5fffffffffffff6f669daff1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c4c51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001650000000000000b0bfbed671c",
    x"0209000000000000025a00000000000000fb335f911c",
    x"030b000000000000025afffffffffffff50003eab51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc0f51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30ea1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd0f291c",
    x"070a0000000000000155fffffffffffff9ef35ece21c",
    x"0802000000000000029afffffffffffff6f669dafc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266c4c11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed681c",
    x"0209000000000000015600000000000000fb335f8b1c",
    x"030b0000000000000156fffffffffffff50003eab61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dc0f31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30e71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd0f231c",
    x"070a00000000000002a9fffffffffffff9ef35ecdf1c",
    x"08020000000000000156fffffffffffff6f669dafa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c4bd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed691c",
    x"0209000000000000031f00000000000000fb335f851c",
    x"030b000000000000031ffffffffffffff50003eab61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc0f01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f30e31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0f1c1c",
    x"070a000000000000031ffffffffffffff9ef35ecdb1c",
    x"0802000000000000031ffffffffffffff6f669daf81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c4b91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed6a1c",
    x"020900000000000000ae00000000000000fb335f801c",
    x"030b00000000000000aefffffffffffff50003eab71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc0ee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f30e01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0f161c",
    x"070a00000000000000aefffffffffffff9ef35ecd71c",
    x"080200000000000000aefffffffffffff6f669daf51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c4b51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed6b1c",
    x"020900000000000001a400000000000000fb335f7a1c",
    x"030b00000000000001a4fffffffffffff50003eab81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc0eb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f30dc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0f101c",
    x"070a00000000000001a4fffffffffffff9ef35ecd31c",
    x"080200000000000001a4fffffffffffff6f669daf31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266c4b11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbed6c1c",
    x"0209000000000000025a00000000000000fb335f751c",
    x"030b000000000000025afffffffffffff50003eab91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc0e91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f30d91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd0f0a1c",
    x"070a000000000000025afffffffffffff9ef35ecd01c",
    x"0802000000000000025afffffffffffff6f669daf01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4ac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed6d1c",
    x"020900000000000002aa00000000000000fb335f6f1c",
    x"030b00000000000002aafffffffffffff50003eaba1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0e61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30d51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0f041c",
    x"070a00000000000002aafffffffffffff9ef35eccc1c",
    x"080200000000000002aafffffffffffff6f669daee1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c4a81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbed6f1c",
    x"0209000000000000029a00000000000000fb335f691c",
    x"030b000000000000029afffffffffffff50003eabb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc0e41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f30d11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd0efd1c",
    x"070a000000000000029afffffffffffff9ef35ecc81c",
    x"0802000000000000029afffffffffffff6f669daeb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4a41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed701c",
    x"020900000000000002aa00000000000000fb335f641c",
    x"030b00000000000002aafffffffffffff50003eabc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0e11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30ce1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ef71c",
    x"070a00000000000002aafffffffffffff9ef35ecc41c",
    x"080200000000000002aafffffffffffff6f669dae91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4a01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed711c",
    x"020900000000000002aa00000000000000fb335f5e1c",
    x"030b00000000000002aafffffffffffff50003eabd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0de1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30ca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ef11c",
    x"070a00000000000002aafffffffffffff9ef35ecc11c",
    x"080200000000000002aafffffffffffff6f669dae71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c49c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed721c",
    x"020900000000000002aa00000000000000fb335f581c",
    x"030b00000000000002aafffffffffffff50003eabd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0dc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30c71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0eeb1c",
    x"070a00000000000002aafffffffffffff9ef35ecbd1c",
    x"080200000000000002aafffffffffffff6f669dae41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4981c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed731c",
    x"020900000000000002aa00000000000000fb335f531c",
    x"030b00000000000002aafffffffffffff50003eabe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0d91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30c31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ee51c",
    x"070a00000000000002aafffffffffffff9ef35ecb91c",
    x"080200000000000002aafffffffffffff6f669dae21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed741c",
    x"020900000000000002aa00000000000000fb335f4d1c",
    x"030b00000000000002aafffffffffffff50003eabf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0d71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30bf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ede1c",
    x"070a00000000000002aafffffffffffff9ef35ecb51c",
    x"080200000000000002aafffffffffffff6f669dadf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c48f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed751c",
    x"020900000000000002aa00000000000000fb335f481c",
    x"030b00000000000002aafffffffffffff50003eac01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0d41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30bc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ed81c",
    x"070a00000000000002aafffffffffffff9ef35ecb21c",
    x"080200000000000002aafffffffffffff6f669dadd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c48b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed771c",
    x"020900000000000002aa00000000000000fb335f421c",
    x"030b00000000000002aafffffffffffff50003eac11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0d21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30b81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ed21c",
    x"070a00000000000002aafffffffffffff9ef35ecae1c",
    x"080200000000000002aafffffffffffff6f669dadb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266c4871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbed781c",
    x"0209000000000000016600000000000000fb335f3c1c",
    x"030b0000000000000166fffffffffffff50003eac21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dc0cf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f30b51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd0ecc1c",
    x"070a0000000000000166fffffffffffff9ef35ecaa1c",
    x"08020000000000000166fffffffffffff6f669dad81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed791c",
    x"0209000000000000015500000000000000fb335f371c",
    x"030b0000000000000155fffffffffffff50003eac31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0cd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30b11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ec61c",
    x"070a0000000000000155fffffffffffff9ef35eca61c",
    x"08020000000000000155fffffffffffff6f669dad61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c47f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed7a1c",
    x"0209000000000000015500000000000000fb335f311c",
    x"030b0000000000000155fffffffffffff50003eac41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0ca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30ad1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ebf1c",
    x"070a0000000000000155fffffffffffff9ef35eca31c",
    x"08020000000000000155fffffffffffff6f669dad31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c47b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed7b1c",
    x"0209000000000000015500000000000000fb335f2b1c",
    x"030b0000000000000155fffffffffffff50003eac41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0c81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30aa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0eb91c",
    x"070a0000000000000155fffffffffffff9ef35ec9f1c",
    x"08020000000000000155fffffffffffff6f669dad11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed7c1c",
    x"0209000000000000015500000000000000fb335f261c",
    x"030b0000000000000155fffffffffffff50003eac51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0c51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30a61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0eb31c",
    x"070a0000000000000155fffffffffffff9ef35ec9b1c",
    x"08020000000000000155fffffffffffff6f669dace1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed7d1c",
    x"0209000000000000015500000000000000fb335f201c",
    x"030b0000000000000155fffffffffffff50003eac61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0c31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30a31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ead1c",
    x"070a0000000000000155fffffffffffff9ef35ec971c",
    x"08020000000000000155fffffffffffff6f669dacc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c46e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbed7f1c",
    x"0209000000000000015900000000000000fb335f1b1c",
    x"030b0000000000000159fffffffffffff50003eac71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dc0c01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f309f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd0ea71c",
    x"070a0000000000000159fffffffffffff9ef35ec941c",
    x"08020000000000000159fffffffffffff6f669daca1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c46a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed801c",
    x"0209000000000000031f00000000000000fb335f151c",
    x"030b000000000000031ffffffffffffff50003eac81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc0bd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f309c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0ea11c",
    x"070a000000000000031ffffffffffffff9ef35ec901c",
    x"0802000000000000031ffffffffffffff6f669dac71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c4661c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed811c",
    x"020900000000000000ae00000000000000fb335f0f1c",
    x"030b00000000000000aefffffffffffff50003eac91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc0bb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f30981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0e9a1c",
    x"070a00000000000000aefffffffffffff9ef35ec8c1c",
    x"080200000000000000aefffffffffffff6f669dac51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c4621c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed821c",
    x"020900000000000001a400000000000000fb335f0a1c",
    x"030b00000000000001a4fffffffffffff50003eaca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc0b81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f30941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0e941c",
    x"070a00000000000001a4fffffffffffff9ef35ec891c",
    x"080200000000000001a4fffffffffffff6f669dac21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c45d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbed831c",
    x"0209000000000000029a00000000000000fb335f041c",
    x"030b000000000000029afffffffffffff50003eaca1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc0b61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f30911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd0e8e1c",
    x"070a000000000000029afffffffffffff9ef35ec851c",
    x"0802000000000000029afffffffffffff6f669dac01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c4591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbed841c",
    x"0209000000000000016a00000000000000fb335efe1c",
    x"030b000000000000016afffffffffffff50003eacb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dc0b31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f308d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd0e881c",
    x"070a000000000000016afffffffffffff9ef35ec811c",
    x"0802000000000000016afffffffffffff6f669dabd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed851c",
    x"020900000000000002aa00000000000000fb335ef91c",
    x"030b00000000000002aafffffffffffff50003eacc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0b11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f308a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e821c",
    x"070a00000000000002aafffffffffffff9ef35ec7d1c",
    x"080200000000000002aafffffffffffff6f669dabb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed871c",
    x"020900000000000002aa00000000000000fb335ef31c",
    x"030b00000000000002aafffffffffffff50003eacd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0ae1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e7b1c",
    x"070a00000000000002aafffffffffffff9ef35ec7a1c",
    x"080200000000000002aafffffffffffff6f669dab91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c44d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed881c",
    x"020900000000000002aa00000000000000fb335eee1c",
    x"030b00000000000002aafffffffffffff50003eace1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0ac1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e751c",
    x"070a00000000000002aafffffffffffff9ef35ec761c",
    x"080200000000000002aafffffffffffff6f669dab61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4491c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed891c",
    x"020900000000000002aa00000000000000fb335ee81c",
    x"030b00000000000002aafffffffffffff50003eacf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0a91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f307f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e6f1c",
    x"070a00000000000002aafffffffffffff9ef35ec721c",
    x"080200000000000002aafffffffffffff6f669dab41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed8a1c",
    x"020900000000000002aa00000000000000fb335ee21c",
    x"030b00000000000002aafffffffffffff50003ead01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0a71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f307b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e691c",
    x"070a00000000000002aafffffffffffff9ef35ec6e1c",
    x"080200000000000002aafffffffffffff6f669dab11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed8b1c",
    x"020900000000000002aa00000000000000fb335edd1c",
    x"030b00000000000002aafffffffffffff50003ead11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0a41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e631c",
    x"070a00000000000002aafffffffffffff9ef35ec6b1c",
    x"080200000000000002aafffffffffffff6f669daaf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c43c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed8c1c",
    x"020900000000000002aa00000000000000fb335ed71c",
    x"030b00000000000002aafffffffffffff50003ead11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0a21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e5c1c",
    x"070a00000000000002aafffffffffffff9ef35ec671c",
    x"080200000000000002aafffffffffffff6f669daac1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed8d1c",
    x"020900000000000002aa00000000000000fb335ed21c",
    x"030b00000000000002aafffffffffffff50003ead21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc09f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30711c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e561c",
    x"070a00000000000002aafffffffffffff9ef35ec631c",
    x"080200000000000002aafffffffffffff6f669daaa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed8f1c",
    x"020900000000000002aa00000000000000fb335ecc1c",
    x"030b00000000000002aafffffffffffff50003ead31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc09d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f306d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e501c",
    x"070a00000000000002aafffffffffffff9ef35ec5f1c",
    x"080200000000000002aafffffffffffff6f669daa81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed901c",
    x"020900000000000002aa00000000000000fb335ec61c",
    x"030b00000000000002aafffffffffffff50003ead41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc09a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e4a1c",
    x"070a00000000000002aafffffffffffff9ef35ec5c1c",
    x"080200000000000002aafffffffffffff6f669daa51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c42c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed911c",
    x"020900000000000002aa00000000000000fb335ec11c",
    x"030b00000000000002aafffffffffffff50003ead51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e441c",
    x"070a00000000000002aafffffffffffff9ef35ec581c",
    x"080200000000000002aafffffffffffff6f669daa31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed921c",
    x"020900000000000002aa00000000000000fb335ebb1c",
    x"030b00000000000002aafffffffffffff50003ead61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0951c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f30621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e3e1c",
    x"070a00000000000002aafffffffffffff9ef35ec541c",
    x"080200000000000002aafffffffffffff6f669daa01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c4231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbed931c",
    x"020900000000000002aa00000000000000fb335eb51c",
    x"030b00000000000002aafffffffffffff50003ead71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0921c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f305f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0e371c",
    x"070a00000000000002aafffffffffffff9ef35ec501c",
    x"080200000000000002aafffffffffffff6f669da9e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000025affffffffffffff0266c41f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000025a0000000000000b0bfbed941c",
    x"0209000000000000025a00000000000000fb335eb01c",
    x"030b000000000000025afffffffffffff50003ead81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000025afffffffffffff4099dc0901c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000025a0000000000000b072f305b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000025a0000000000000004cd0e311c",
    x"070a000000000000025afffffffffffff9ef35ec4d1c",
    x"0802000000000000025afffffffffffff6f669da9c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c41b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed951c",
    x"0209000000000000015500000000000000fb335eaa1c",
    x"030b0000000000000155fffffffffffff50003ead81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc08d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0e2b1c",
    x"070a0000000000000155fffffffffffff9ef35ec491c",
    x"08020000000000000155fffffffffffff6f669da991c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c4171c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbed971c",
    x"0209000000000000031f00000000000000fb335ea51c",
    x"030b000000000000031ffffffffffffff50003ead91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc08b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f30541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0e251c",
    x"070a000000000000031ffffffffffffff9ef35ec451c",
    x"0802000000000000031ffffffffffffff6f669da971c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c4131c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbed981c",
    x"020900000000000000ae00000000000000fb335e9f1c",
    x"030b00000000000000aefffffffffffff50003eada1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc0881c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f30501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0e1f1c",
    x"070a00000000000000aefffffffffffff9ef35ec411c",
    x"080200000000000000aefffffffffffff6f669da941c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c40e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbed991c",
    x"020900000000000001a400000000000000fb335e991c",
    x"030b00000000000001a4fffffffffffff50003eadb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc0861c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f304d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0e181c",
    x"070a00000000000001a4fffffffffffff9ef35ec3e1c",
    x"080200000000000001a4fffffffffffff6f669da921c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000019affffffffffffff0266c40a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000019a0000000000000b0bfbed9a1c",
    x"0209000000000000019a00000000000000fb335e941c",
    x"030b000000000000019afffffffffffff50003eadc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000019afffffffffffff4099dc0831c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000019a0000000000000b072f30491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000019a0000000000000004cd0e121c",
    x"070a000000000000019afffffffffffff9ef35ec3a1c",
    x"0802000000000000019afffffffffffff6f669da8f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4061c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed9b1c",
    x"0209000000000000015500000000000000fb335e8e1c",
    x"030b0000000000000155fffffffffffff50003eadd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0811c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30451c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0e0c1c",
    x"070a0000000000000155fffffffffffff9ef35ec361c",
    x"08020000000000000155fffffffffffff6f669da8d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c4021c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed9c1c",
    x"0209000000000000015500000000000000fb335e881c",
    x"030b0000000000000155fffffffffffff50003eade1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc07e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0e061c",
    x"070a0000000000000155fffffffffffff9ef35ec321c",
    x"08020000000000000155fffffffffffff6f669da8b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3fe1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed9d1c",
    x"0209000000000000015500000000000000fb335e831c",
    x"030b0000000000000155fffffffffffff50003eade1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc07c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f303e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0e001c",
    x"070a0000000000000155fffffffffffff9ef35ec2f1c",
    x"08020000000000000155fffffffffffff6f669da881c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3fa1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbed9f1c",
    x"0209000000000000015500000000000000fb335e7d1c",
    x"030b0000000000000155fffffffffffff50003eadf1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0791c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f303b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0df91c",
    x"070a0000000000000155fffffffffffff9ef35ec2b1c",
    x"08020000000000000155fffffffffffff6f669da861c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3f61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda01c",
    x"0209000000000000015500000000000000fb335e781c",
    x"030b0000000000000155fffffffffffff50003eae01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0761c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0df31c",
    x"070a0000000000000155fffffffffffff9ef35ec271c",
    x"08020000000000000155fffffffffffff6f669da831c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3f11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda11c",
    x"0209000000000000015500000000000000fb335e721c",
    x"030b0000000000000155fffffffffffff50003eae11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0741c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ded1c",
    x"070a0000000000000155fffffffffffff9ef35ec231c",
    x"08020000000000000155fffffffffffff6f669da811c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3ed1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda21c",
    x"0209000000000000015500000000000000fb335e6c1c",
    x"030b0000000000000155fffffffffffff50003eae21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0711c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30301c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0de71c",
    x"070a0000000000000155fffffffffffff9ef35ec201c",
    x"08020000000000000155fffffffffffff6f669da7e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3e91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda31c",
    x"0209000000000000015500000000000000fb335e671c",
    x"030b0000000000000155fffffffffffff50003eae31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc06f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f302c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0de11c",
    x"070a0000000000000155fffffffffffff9ef35ec1c1c",
    x"08020000000000000155fffffffffffff6f669da7c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3e51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda41c",
    x"0209000000000000015500000000000000fb335e611c",
    x"030b0000000000000155fffffffffffff50003eae41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc06c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0dda1c",
    x"070a0000000000000155fffffffffffff9ef35ec181c",
    x"08020000000000000155fffffffffffff6f669da7a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3e11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda51c",
    x"0209000000000000015500000000000000fb335e5b1c",
    x"030b0000000000000155fffffffffffff50003eae51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc06a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30251c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0dd41c",
    x"070a0000000000000155fffffffffffff9ef35ec141c",
    x"08020000000000000155fffffffffffff6f669da771c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3dd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda71c",
    x"0209000000000000015500000000000000fb335e561c",
    x"030b0000000000000155fffffffffffff50003eae51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0671c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30221c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0dce1c",
    x"070a0000000000000155fffffffffffff9ef35ec111c",
    x"08020000000000000155fffffffffffff6f669da751c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3d81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda81c",
    x"0209000000000000015500000000000000fb335e501c",
    x"030b0000000000000155fffffffffffff50003eae61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0651c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f301e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0dc81c",
    x"070a0000000000000155fffffffffffff9ef35ec0d1c",
    x"08020000000000000155fffffffffffff6f669da721c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3d41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbeda91c",
    x"0209000000000000015500000000000000fb335e4b1c",
    x"030b0000000000000155fffffffffffff50003eae71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0621c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f301a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0dc21c",
    x"070a0000000000000155fffffffffffff9ef35ec091c",
    x"08020000000000000155fffffffffffff6f669da701c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3d01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedaa1c",
    x"0209000000000000015500000000000000fb335e451c",
    x"030b0000000000000155fffffffffffff50003eae81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0601c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0dbc1c",
    x"070a0000000000000155fffffffffffff9ef35ec051c",
    x"08020000000000000155fffffffffffff6f669da6d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3cc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedab1c",
    x"0209000000000000015500000000000000fb335e3f1c",
    x"030b0000000000000155fffffffffffff50003eae91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc05d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30131c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0db51c",
    x"070a0000000000000155fffffffffffff9ef35ec021c",
    x"08020000000000000155fffffffffffff6f669da6b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3c81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedac1c",
    x"0209000000000000015500000000000000fb335e3a1c",
    x"030b0000000000000155fffffffffffff50003eaea1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc05a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f30101c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0daf1c",
    x"070a0000000000000155fffffffffffff9ef35ebfe1c",
    x"08020000000000000155fffffffffffff6f669da691c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c3c41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbedad1c",
    x"0209000000000000031f00000000000000fb335e341c",
    x"030b000000000000031ffffffffffffff50003eaeb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc0581c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f300c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0da91c",
    x"070a000000000000031ffffffffffffff9ef35ebfa1c",
    x"0802000000000000031ffffffffffffff6f669da661c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c3c01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbedaf1c",
    x"020900000000000000ae00000000000000fb335e2f1c",
    x"030b00000000000000aefffffffffffff50003eaeb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc0551c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f30091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0da31c",
    x"070a00000000000000aefffffffffffff9ef35ebf71c",
    x"080200000000000000aefffffffffffff6f669da641c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c3bb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbedb01c",
    x"020900000000000001a400000000000000fb335e291c",
    x"030b00000000000001a4fffffffffffff50003eaec1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc0531c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f30051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0d9d1c",
    x"070a00000000000001a4fffffffffffff9ef35ebf31c",
    x"080200000000000001a4fffffffffffff6f669da611c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000156ffffffffffffff0266c3b71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001560000000000000b0bfbedb11c",
    x"0209000000000000015600000000000000fb335e231c",
    x"030b0000000000000156fffffffffffff50003eaed1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000156fffffffffffff4099dc0501c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001560000000000000b072f30011c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001560000000000000004cd0d961c",
    x"070a0000000000000156fffffffffffff9ef35ebef1c",
    x"08020000000000000156fffffffffffff6f669da5f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3b31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedb21c",
    x"0209000000000000015500000000000000fb335e1e1c",
    x"030b0000000000000155fffffffffffff50003eaee1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc04e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ffe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0d901c",
    x"070a0000000000000155fffffffffffff9ef35ebeb1c",
    x"08020000000000000155fffffffffffff6f669da5c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c3af1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbedb31c",
    x"0209000000000000029a00000000000000fb335e181c",
    x"030b000000000000029afffffffffffff50003eaef1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dc04b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f2ffa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd0d8a1c",
    x"070a000000000000029afffffffffffff9ef35ebe81c",
    x"0802000000000000029afffffffffffff6f669da5a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3ab1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedb41c",
    x"020900000000000002aa00000000000000fb335e121c",
    x"030b00000000000002aafffffffffffff50003eaf01c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0491c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2ff71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d841c",
    x"070a00000000000002aafffffffffffff9ef35ebe41c",
    x"080200000000000002aafffffffffffff6f669da581c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3a71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedb51c",
    x"020900000000000002aa00000000000000fb335e0d1c",
    x"030b00000000000002aafffffffffffff50003eaf11c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0461c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2ff31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d7e1c",
    x"070a00000000000002aafffffffffffff9ef35ebe01c",
    x"080200000000000002aafffffffffffff6f669da551c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3a21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedb71c",
    x"020900000000000002aa00000000000000fb335e071c",
    x"030b00000000000002aafffffffffffff50003eaf21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0441c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fef1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d771c",
    x"070a00000000000002aafffffffffffff9ef35ebdc1c",
    x"080200000000000002aafffffffffffff6f669da531c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c39e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedb81c",
    x"020900000000000002aa00000000000000fb335e021c",
    x"030b00000000000002aafffffffffffff50003eaf21c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0411c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d711c",
    x"070a00000000000002aafffffffffffff9ef35ebd91c",
    x"080200000000000002aafffffffffffff6f669da501c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c39a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedb91c",
    x"020900000000000002aa00000000000000fb335dfc1c",
    x"030b00000000000002aafffffffffffff50003eaf31c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc03f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fe81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d6b1c",
    x"070a00000000000002aafffffffffffff9ef35ebd51c",
    x"080200000000000002aafffffffffffff6f669da4e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3961c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedba1c",
    x"020900000000000002aa00000000000000fb335df61c",
    x"030b00000000000002aafffffffffffff50003eaf41c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc03c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fe51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d651c",
    x"070a00000000000002aafffffffffffff9ef35ebd11c",
    x"080200000000000002aafffffffffffff6f669da4b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3921c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedbb1c",
    x"020900000000000002aa00000000000000fb335df11c",
    x"030b00000000000002aafffffffffffff50003eaf51c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0391c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fe11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d5f1c",
    x"070a00000000000002aafffffffffffff9ef35ebcd1c",
    x"080200000000000002aafffffffffffff6f669da491c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c38e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedbc1c",
    x"020900000000000002aa00000000000000fb335deb1c",
    x"030b00000000000002aafffffffffffff50003eaf61c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0371c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fde1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d581c",
    x"070a00000000000002aafffffffffffff9ef35ebca1c",
    x"080200000000000002aafffffffffffff6f669da471c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c38a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedbd1c",
    x"020900000000000002aa00000000000000fb335de51c",
    x"030b00000000000002aafffffffffffff50003eaf71c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0341c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fda1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d521c",
    x"070a00000000000002aafffffffffffff9ef35ebc61c",
    x"080200000000000002aafffffffffffff6f669da441c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3851c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedbf1c",
    x"020900000000000002aa00000000000000fb335de01c",
    x"030b00000000000002aafffffffffffff50003eaf81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0321c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fd61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d4c1c",
    x"070a00000000000002aafffffffffffff9ef35ebc21c",
    x"080200000000000002aafffffffffffff6f669da421c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3811c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedc01c",
    x"020900000000000002aa00000000000000fb335dda1c",
    x"030b00000000000002aafffffffffffff50003eaf81c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc02f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fd31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d461c",
    x"070a00000000000002aafffffffffffff9ef35ebbe1c",
    x"080200000000000002aafffffffffffff6f669da3f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c37d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedc11c",
    x"020900000000000002aa00000000000000fb335dd51c",
    x"030b00000000000002aafffffffffffff50003eaf91c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc02d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fcf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d401c",
    x"070a00000000000002aafffffffffffff9ef35ebbb1c",
    x"080200000000000002aafffffffffffff6f669da3d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000026affffffffffffff0266c3791c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000026a0000000000000b0bfbedc21c",
    x"0209000000000000026a00000000000000fb335dcf1c",
    x"030b000000000000026afffffffffffff50003eafa1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000026afffffffffffff4099dc02a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000026a0000000000000b072f2fcc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000026a0000000000000004cd0d391c",
    x"070a000000000000026afffffffffffff9ef35ebb71c",
    x"0802000000000000026afffffffffffff6f669da3b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c3751c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedc31c",
    x"0209000000000000015500000000000000fb335dc91c",
    x"030b0000000000000155fffffffffffff50003eafb1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dc0281c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2fc81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0d331c",
    x"070a0000000000000155fffffffffffff9ef35ebb31c",
    x"08020000000000000155fffffffffffff6f669da381c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c3711c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbedc41c",
    x"0209000000000000031f00000000000000fb335dc41c",
    x"030b000000000000031ffffffffffffff50003eafc1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dc0251c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2fc41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0d2d1c",
    x"070a000000000000031ffffffffffffff9ef35ebaf1c",
    x"0802000000000000031ffffffffffffff6f669da361c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c36c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbedc61c",
    x"020900000000000000ae00000000000000fb335dbe1c",
    x"030b00000000000000aefffffffffffff50003eafd1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dc0231c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2fc11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0d271c",
    x"070a00000000000000aefffffffffffff9ef35ebac1c",
    x"080200000000000000aefffffffffffff6f669da331c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c3681c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbedc71c",
    x"020900000000000001a400000000000000fb335db81c",
    x"030b00000000000001a4fffffffffffff50003eafe1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dc0201c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2fbd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0d211c",
    x"070a00000000000001a4fffffffffffff9ef35eba81c",
    x"080200000000000001a4fffffffffffff6f669da311c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000256ffffffffffffff0266c3641c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002560000000000000b0bfbedc81c",
    x"0209000000000000025600000000000000fb335db31c",
    x"030b0000000000000256fffffffffffff50003eaff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000256fffffffffffff4099dc01d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002560000000000000b072f2fba1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002560000000000000004cd0d1b1c",
    x"070a0000000000000256fffffffffffff9ef35eba41c",
    x"08020000000000000256fffffffffffff6f669da2e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3601c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedc91c",
    x"020900000000000002aa00000000000000fb335dad1c",
    x"030b00000000000002aafffffffffffff50003eaff1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc01b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fb61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d141c",
    x"070a00000000000002aafffffffffffff9ef35eba01c",
    x"080200000000000002aafffffffffffff6f669da2c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c35c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedca1c",
    x"020900000000000002aa00000000000000fb335da81c",
    x"030b00000000000002aafffffffffffff50003eb001c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0181c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fb31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d0e1c",
    x"070a00000000000002aafffffffffffff9ef35eb9d1c",
    x"080200000000000002aafffffffffffff6f669da2a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3581c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedcb1c",
    x"020900000000000002aa00000000000000fb335da21c",
    x"030b00000000000002aafffffffffffff50003eb011c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0161c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2faf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d081c",
    x"070a00000000000002aafffffffffffff9ef35eb991c",
    x"080200000000000002aafffffffffffff6f669da271c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3541c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedcc1c",
    x"020900000000000002aa00000000000000fb335d9c1c",
    x"030b00000000000002aafffffffffffff50003eb021c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0131c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fab1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0d021c",
    x"070a00000000000002aafffffffffffff9ef35eb951c",
    x"080200000000000002aafffffffffffff6f669da251c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c34f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedce1c",
    x"020900000000000002aa00000000000000fb335d971c",
    x"030b00000000000002aafffffffffffff50003eb031c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0111c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fa81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cfc1c",
    x"070a00000000000002aafffffffffffff9ef35eb911c",
    x"080200000000000002aafffffffffffff6f669da221c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c34b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedcf1c",
    x"020900000000000002aa00000000000000fb335d911c",
    x"030b00000000000002aafffffffffffff50003eb041c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc00e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fa41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cf51c",
    x"070a00000000000002aafffffffffffff9ef35eb8e1c",
    x"080200000000000002aafffffffffffff6f669da201c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3471c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd01c",
    x"020900000000000002aa00000000000000fb335d8b1c",
    x"030b00000000000002aafffffffffffff50003eb051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc00c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2fa11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cef1c",
    x"070a00000000000002aafffffffffffff9ef35eb8a1c",
    x"080200000000000002aafffffffffffff6f669da1d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3431c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd11c",
    x"020900000000000002aa00000000000000fb335d861c",
    x"030b00000000000002aafffffffffffff50003eb051c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0091c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f9d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ce91c",
    x"070a00000000000002aafffffffffffff9ef35eb861c",
    x"080200000000000002aafffffffffffff6f669da1b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c33f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd21c",
    x"020900000000000002aa00000000000000fb335d801c",
    x"030b00000000000002aafffffffffffff50003eb061c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0071c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f991c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ce31c",
    x"070a00000000000002aafffffffffffff9ef35eb821c",
    x"080200000000000002aafffffffffffff6f669da191c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c33b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd31c",
    x"020900000000000002aa00000000000000fb335d7b1c",
    x"030b00000000000002aafffffffffffff50003eb071c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0041c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f961c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cdd1c",
    x"070a00000000000002aafffffffffffff9ef35eb7f1c",
    x"080200000000000002aafffffffffffff6f669da161c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3361c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd41c",
    x"020900000000000002aa00000000000000fb335d751c",
    x"030b00000000000002aafffffffffffff50003eb081c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dc0021c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f921c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cd61c",
    x"070a00000000000002aafffffffffffff9ef35eb7b1c",
    x"080200000000000002aafffffffffffff6f669da141c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3321c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd61c",
    x"020900000000000002aa00000000000000fb335d6f1c",
    x"030b00000000000002aafffffffffffff50003eb091c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfff1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f8f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cd01c",
    x"070a00000000000002aafffffffffffff9ef35eb771c",
    x"080200000000000002aafffffffffffff6f669da111c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c32e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd71c",
    x"020900000000000002aa00000000000000fb335d6a1c",
    x"030b00000000000002aafffffffffffff50003eb0a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbffc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f8b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cca1c",
    x"070a00000000000002aafffffffffffff9ef35eb731c",
    x"080200000000000002aafffffffffffff6f669da0f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c32a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedd81c",
    x"020900000000000002aa00000000000000fb335d641c",
    x"030b00000000000002aafffffffffffff50003eb0b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbffa1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f881c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cc41c",
    x"070a00000000000002aafffffffffffff9ef35eb701c",
    x"080200000000000002aafffffffffffff6f669da0c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000029affffffffffffff0266c3261c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000029a0000000000000b0bfbedd91c",
    x"0209000000000000029a00000000000000fb335d5e1c",
    x"030b000000000000029afffffffffffff50003eb0b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000029afffffffffffff4099dbff71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000029a0000000000000b072f2f841c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000029a0000000000000004cd0cbe1c",
    x"070a000000000000029afffffffffffff9ef35eb6c1c",
    x"0802000000000000029afffffffffffff6f669da0a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3221c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedda1c",
    x"020900000000000002aa00000000000000fb335d591c",
    x"030b00000000000002aafffffffffffff50003eb0c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbff51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f801c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0cb71c",
    x"070a00000000000002aafffffffffffff9ef35eb681c",
    x"080200000000000002aafffffffffffff6f669da081c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c31e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbeddb1c",
    x"0209000000000000031f00000000000000fb335d531c",
    x"030b000000000000031ffffffffffffff50003eb0d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbff21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2f7d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0cb11c",
    x"070a000000000000031ffffffffffffff9ef35eb641c",
    x"0802000000000000031ffffffffffffff6f669da051c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c3191c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbeddc1c",
    x"020900000000000000ae00000000000000fb335d4e1c",
    x"030b00000000000000aefffffffffffff50003eb0e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbff01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2f791c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0cab1c",
    x"070a00000000000000aefffffffffffff9ef35eb611c",
    x"080200000000000000aefffffffffffff6f669da031c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c3151c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbedde1c",
    x"020900000000000001a400000000000000fb335d481c",
    x"030b00000000000001a4fffffffffffff50003eb0f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbfed1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2f761c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0ca51c",
    x"070a00000000000001a4fffffffffffff9ef35eb5d1c",
    x"080200000000000001a4fffffffffffff6f669da001c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000296ffffffffffffff0266c3111c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002960000000000000b0bfbeddf1c",
    x"0209000000000000029600000000000000fb335d421c",
    x"030b0000000000000296fffffffffffff50003eb101c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000296fffffffffffff4099dbfeb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002960000000000000b072f2f721c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002960000000000000004cd0c9f1c",
    x"070a0000000000000296fffffffffffff9ef35eb591c",
    x"08020000000000000296fffffffffffff6f669d9fe1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c30d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede01c",
    x"020900000000000002aa00000000000000fb335d3d1c",
    x"030b00000000000002aafffffffffffff50003eb111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfe81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f6e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c991c",
    x"070a00000000000002aafffffffffffff9ef35eb551c",
    x"080200000000000002aafffffffffffff6f669d9fb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a9ffffffffffffff0266c3091c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a90000000000000b0bfbede11c",
    x"020900000000000002a900000000000000fb335d371c",
    x"030b00000000000002a9fffffffffffff50003eb111c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a9fffffffffffff4099dbfe61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a90000000000000b072f2f6b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a90000000000000004cd0c921c",
    x"070a00000000000002a9fffffffffffff9ef35eb521c",
    x"080200000000000002a9fffffffffffff6f669d9f91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3051c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede21c",
    x"020900000000000002aa00000000000000fb335d321c",
    x"030b00000000000002aafffffffffffff50003eb121c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfe31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f671c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c8c1c",
    x"070a00000000000002aafffffffffffff9ef35eb4e1c",
    x"080200000000000002aafffffffffffff6f669d9f71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c3001c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede31c",
    x"020900000000000002aa00000000000000fb335d2c1c",
    x"030b00000000000002aafffffffffffff50003eb131c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfe01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f641c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c861c",
    x"070a00000000000002aafffffffffffff9ef35eb4a1c",
    x"080200000000000002aafffffffffffff6f669d9f41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2fc1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede41c",
    x"020900000000000002aa00000000000000fb335d261c",
    x"030b00000000000002aafffffffffffff50003eb141c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfde1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f601c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c801c",
    x"070a00000000000002aafffffffffffff9ef35eb461c",
    x"080200000000000002aafffffffffffff6f669d9f21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2f81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede61c",
    x"020900000000000002aa00000000000000fb335d211c",
    x"030b00000000000002aafffffffffffff50003eb151c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfdb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f5d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c7a1c",
    x"070a00000000000002aafffffffffffff9ef35eb431c",
    x"080200000000000002aafffffffffffff6f669d9ef1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2f41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede71c",
    x"020900000000000002aa00000000000000fb335d1b1c",
    x"030b00000000000002aafffffffffffff50003eb161c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfd91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f591c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c731c",
    x"070a00000000000002aafffffffffffff9ef35eb3f1c",
    x"080200000000000002aafffffffffffff6f669d9ed1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2f01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede81c",
    x"020900000000000002aa00000000000000fb335d151c",
    x"030b00000000000002aafffffffffffff50003eb171c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfd61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f551c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c6d1c",
    x"070a00000000000002aafffffffffffff9ef35eb3b1c",
    x"080200000000000002aafffffffffffff6f669d9ea1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2ec1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbede91c",
    x"020900000000000002aa00000000000000fb335d101c",
    x"030b00000000000002aafffffffffffff50003eb181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfd41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f521c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c671c",
    x"070a00000000000002aafffffffffffff9ef35eb371c",
    x"080200000000000002aafffffffffffff6f669d9e81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2e81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedea1c",
    x"020900000000000002aa00000000000000fb335d0a1c",
    x"030b00000000000002aafffffffffffff50003eb181c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfd11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f4e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c611c",
    x"070a00000000000002aafffffffffffff9ef35eb341c",
    x"080200000000000002aafffffffffffff6f669d9e61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2e31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedeb1c",
    x"020900000000000002aa00000000000000fb335d051c",
    x"030b00000000000002aafffffffffffff50003eb191c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfcf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f4b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c5b1c",
    x"070a00000000000002aafffffffffffff9ef35eb301c",
    x"080200000000000002aafffffffffffff6f669d9e31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2df1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedec1c",
    x"020900000000000002aa00000000000000fb335cff1c",
    x"030b00000000000002aafffffffffffff50003eb1a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfcc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f471c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c541c",
    x"070a00000000000002aafffffffffffff9ef35eb2c1c",
    x"080200000000000002aafffffffffffff6f669d9e11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2db1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedee1c",
    x"020900000000000002aa00000000000000fb335cf91c",
    x"030b00000000000002aafffffffffffff50003eb1b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f441c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c4e1c",
    x"070a00000000000002aafffffffffffff9ef35eb281c",
    x"080200000000000002aafffffffffffff6f669d9de1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c2d71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbedef1c",
    x"020900000000000002aa00000000000000fb335cf41c",
    x"030b00000000000002aafffffffffffff50003eb1c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbfc71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2f401c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0c481c",
    x"070a00000000000002aafffffffffffff9ef35eb251c",
    x"080200000000000002aafffffffffffff6f669d9dc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000015affffffffffffff0266c2d31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000015a0000000000000b0bfbedf01c",
    x"0209000000000000015a00000000000000fb335cee1c",
    x"030b000000000000015afffffffffffff50003eb1d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000015afffffffffffff4099dbfc41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000015a0000000000000b072f2f3c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000015a0000000000000004cd0c421c",
    x"070a000000000000015afffffffffffff9ef35eb211c",
    x"0802000000000000015afffffffffffff6f669d9d91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2cf1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedf11c",
    x"0209000000000000015500000000000000fb335ce81c",
    x"030b0000000000000155fffffffffffff50003eb1e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfc21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f391c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0c3c1c",
    x"070a0000000000000155fffffffffffff9ef35eb1d1c",
    x"08020000000000000155fffffffffffff6f669d9d71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c2ca1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbedf21c",
    x"0209000000000000031f00000000000000fb335ce31c",
    x"030b000000000000031ffffffffffffff50003eb1e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbfbf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2f351c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0c351c",
    x"070a000000000000031ffffffffffffff9ef35eb191c",
    x"0802000000000000031ffffffffffffff6f669d9d51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c2c61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbedf31c",
    x"020900000000000000ae00000000000000fb335cdd1c",
    x"030b00000000000000aefffffffffffff50003eb1f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbfbd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2f321c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0c2f1c",
    x"070a00000000000000aefffffffffffff9ef35eb161c",
    x"080200000000000000aefffffffffffff6f669d9d21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c2c21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbedf41c",
    x"020900000000000001a400000000000000fb335cd81c",
    x"030b00000000000001a4fffffffffffff50003eb201c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbfba1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2f2e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0c291c",
    x"070a00000000000001a4fffffffffffff9ef35eb121c",
    x"080200000000000001a4fffffffffffff6f669d9d01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000196ffffffffffffff0266c2be1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001960000000000000b0bfbedf61c",
    x"0209000000000000019600000000000000fb335cd21c",
    x"030b0000000000000196fffffffffffff50003eb211c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000196fffffffffffff4099dbfb81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001960000000000000b072f2f2a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001960000000000000004cd0c231c",
    x"070a0000000000000196fffffffffffff9ef35eb0e1c",
    x"08020000000000000196fffffffffffff6f669d9cd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2ba1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedf71c",
    x"0209000000000000015500000000000000fb335ccc1c",
    x"030b0000000000000155fffffffffffff50003eb221c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfb51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f271c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0c1d1c",
    x"070a0000000000000155fffffffffffff9ef35eb0a1c",
    x"08020000000000000155fffffffffffff6f669d9cb1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2b61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedf81c",
    x"0209000000000000015500000000000000fb335cc71c",
    x"030b0000000000000155fffffffffffff50003eb231c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfb31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f231c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0c161c",
    x"070a0000000000000155fffffffffffff9ef35eb071c",
    x"08020000000000000155fffffffffffff6f669d9c81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2b21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedf91c",
    x"0209000000000000015500000000000000fb335cc11c",
    x"030b0000000000000155fffffffffffff50003eb241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfb01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f201c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0c101c",
    x"070a0000000000000155fffffffffffff9ef35eb031c",
    x"08020000000000000155fffffffffffff6f669d9c61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2ad1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedfa1c",
    x"0209000000000000015500000000000000fb335cbb1c",
    x"030b0000000000000155fffffffffffff50003eb241c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfad1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f1c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0c0a1c",
    x"070a0000000000000155fffffffffffff9ef35eaff1c",
    x"08020000000000000155fffffffffffff6f669d9c41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2a91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedfb1c",
    x"0209000000000000015500000000000000fb335cb61c",
    x"030b0000000000000155fffffffffffff50003eb251c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfab1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f191c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0c041c",
    x"070a0000000000000155fffffffffffff9ef35eafb1c",
    x"08020000000000000155fffffffffffff6f669d9c11c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2a51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedfd1c",
    x"0209000000000000015500000000000000fb335cb01c",
    x"030b0000000000000155fffffffffffff50003eb261c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfa81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f151c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bfe1c",
    x"070a0000000000000155fffffffffffff9ef35eaf81c",
    x"08020000000000000155fffffffffffff6f669d9bf1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2a11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedfe1c",
    x"0209000000000000015500000000000000fb335cab1c",
    x"030b0000000000000155fffffffffffff50003eb271c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfa61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f111c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bf81c",
    x"070a0000000000000155fffffffffffff9ef35eaf41c",
    x"08020000000000000155fffffffffffff6f669d9bc1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c29d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbedff1c",
    x"0209000000000000015500000000000000fb335ca51c",
    x"030b0000000000000155fffffffffffff50003eb281c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfa31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f0e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bf11c",
    x"070a0000000000000155fffffffffffff9ef35eaf01c",
    x"08020000000000000155fffffffffffff6f669d9ba1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2991c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee001c",
    x"0209000000000000015500000000000000fb335c9f1c",
    x"030b0000000000000155fffffffffffff50003eb291c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbfa11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f0a1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0beb1c",
    x"070a0000000000000155fffffffffffff9ef35eaec1c",
    x"08020000000000000155fffffffffffff6f669d9b71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2951c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee011c",
    x"0209000000000000015500000000000000fb335c9a1c",
    x"030b0000000000000155fffffffffffff50003eb2a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf9e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f071c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0be51c",
    x"070a0000000000000155fffffffffffff9ef35eae91c",
    x"08020000000000000155fffffffffffff6f669d9b51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2901c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee021c",
    x"0209000000000000015500000000000000fb335c941c",
    x"030b0000000000000155fffffffffffff50003eb2a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf9c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f031c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bdf1c",
    x"070a0000000000000155fffffffffffff9ef35eae51c",
    x"08020000000000000155fffffffffffff6f669d9b31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c28c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee031c",
    x"0209000000000000015500000000000000fb335c8e1c",
    x"030b0000000000000155fffffffffffff50003eb2b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf991c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2f001c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bd91c",
    x"070a0000000000000155fffffffffffff9ef35eae11c",
    x"08020000000000000155fffffffffffff6f669d9b01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2881c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee051c",
    x"0209000000000000015500000000000000fb335c891c",
    x"030b0000000000000155fffffffffffff50003eb2c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf971c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2efc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bd21c",
    x"070a0000000000000155fffffffffffff9ef35eadd1c",
    x"08020000000000000155fffffffffffff6f669d9ae1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2841c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee061c",
    x"0209000000000000015500000000000000fb335c831c",
    x"030b0000000000000155fffffffffffff50003eb2d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf941c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ef81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0bcc1c",
    x"070a0000000000000155fffffffffffff9ef35eada1c",
    x"08020000000000000155fffffffffffff6f669d9ab1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a5ffffffffffffff0266c2801c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a50000000000000b0bfbee071c",
    x"020900000000000002a500000000000000fb335c7e1c",
    x"030b00000000000002a5fffffffffffff50003eb2e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a5fffffffffffff4099dbf911c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a50000000000000b072f2ef51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a50000000000000004cd0bc61c",
    x"070a00000000000002a5fffffffffffff9ef35ead61c",
    x"080200000000000002a5fffffffffffff6f669d9a91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c27c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee081c",
    x"020900000000000002aa00000000000000fb335c781c",
    x"030b00000000000002aafffffffffffff50003eb2f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbf8f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2ef11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0bc01c",
    x"070a00000000000002aafffffffffffff9ef35ead21c",
    x"080200000000000002aafffffffffffff6f669d9a61c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c2771c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbee091c",
    x"0209000000000000031f00000000000000fb335c721c",
    x"030b000000000000031ffffffffffffff50003eb301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbf8c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2eee1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0bba1c",
    x"070a000000000000031ffffffffffffff9ef35eace1c",
    x"0802000000000000031ffffffffffffff6f669d9a41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c2731c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbee0a1c",
    x"020900000000000000ae00000000000000fb335c6d1c",
    x"030b00000000000000aefffffffffffff50003eb301c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbf8a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2eea1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0bb31c",
    x"070a00000000000000aefffffffffffff9ef35eacb1c",
    x"080200000000000000aefffffffffffff6f669d9a21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c26f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbee0b1c",
    x"020900000000000001a400000000000000fb335c671c",
    x"030b00000000000001a4fffffffffffff50003eb311c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbf871c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2ee61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0bad1c",
    x"070a00000000000001a4fffffffffffff9ef35eac71c",
    x"080200000000000001a4fffffffffffff6f669d99f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002a6ffffffffffffff0266c26b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002a60000000000000b0bfbee0d1c",
    x"020900000000000002a600000000000000fb335c611c",
    x"030b00000000000002a6fffffffffffff50003eb321c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002a6fffffffffffff4099dbf851c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002a60000000000000b072f2ee31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002a60000000000000004cd0ba71c",
    x"070a00000000000002a6fffffffffffff9ef35eac31c",
    x"080200000000000002a6fffffffffffff6f669d99d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000016affffffffffffff0266c2671c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000016a0000000000000b0bfbee0e1c",
    x"0209000000000000016a00000000000000fb335c5c1c",
    x"030b000000000000016afffffffffffff50003eb331c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000016afffffffffffff4099dbf821c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000016a0000000000000b072f2edf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000016a0000000000000004cd0ba11c",
    x"070a000000000000016afffffffffffff9ef35eabf1c",
    x"0802000000000000016afffffffffffff6f669d99a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000169ffffffffffffff0266c2631c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001690000000000000b0bfbee0f1c",
    x"0209000000000000016900000000000000fb335c561c",
    x"030b0000000000000169fffffffffffff50003eb341c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000169fffffffffffff4099dbf801c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001690000000000000b072f2edc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001690000000000000004cd0b9b1c",
    x"070a0000000000000169fffffffffffff9ef35eabc1c",
    x"08020000000000000169fffffffffffff6f669d9981c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c25f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee101c",
    x"0209000000000000015500000000000000fb335c511c",
    x"030b0000000000000155fffffffffffff50003eb351c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf7d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ed81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b941c",
    x"070a0000000000000155fffffffffffff9ef35eab81c",
    x"08020000000000000155fffffffffffff6f669d9961c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c25a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee111c",
    x"0209000000000000015500000000000000fb335c4b1c",
    x"030b0000000000000155fffffffffffff50003eb361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf7b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ed51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b8e1c",
    x"070a0000000000000155fffffffffffff9ef35eab41c",
    x"08020000000000000155fffffffffffff6f669d9931c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2561c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee121c",
    x"0209000000000000015500000000000000fb335c451c",
    x"030b0000000000000155fffffffffffff50003eb361c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf781c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ed11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b881c",
    x"070a0000000000000155fffffffffffff9ef35eab01c",
    x"08020000000000000155fffffffffffff6f669d9911c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2521c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee131c",
    x"0209000000000000015500000000000000fb335c401c",
    x"030b0000000000000155fffffffffffff50003eb371c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf751c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ecd1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b821c",
    x"070a0000000000000155fffffffffffff9ef35eaad1c",
    x"08020000000000000155fffffffffffff6f669d98e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c24e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee151c",
    x"0209000000000000015500000000000000fb335c3a1c",
    x"030b0000000000000155fffffffffffff50003eb381c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf731c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2eca1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b7c1c",
    x"070a0000000000000155fffffffffffff9ef35eaa91c",
    x"08020000000000000155fffffffffffff6f669d98c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c24a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee161c",
    x"0209000000000000015500000000000000fb335c341c",
    x"030b0000000000000155fffffffffffff50003eb391c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf701c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ec61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b751c",
    x"070a0000000000000155fffffffffffff9ef35eaa51c",
    x"08020000000000000155fffffffffffff6f669d9891c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2461c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee171c",
    x"0209000000000000015500000000000000fb335c2f1c",
    x"030b0000000000000155fffffffffffff50003eb3a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf6e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ec31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b6f1c",
    x"070a0000000000000155fffffffffffff9ef35eaa11c",
    x"08020000000000000155fffffffffffff6f669d9871c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2411c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee181c",
    x"0209000000000000015500000000000000fb335c291c",
    x"030b0000000000000155fffffffffffff50003eb3b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf6b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ebf1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b691c",
    x"070a0000000000000155fffffffffffff9ef35ea9d1c",
    x"08020000000000000155fffffffffffff6f669d9851c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c23d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee191c",
    x"0209000000000000015500000000000000fb335c241c",
    x"030b0000000000000155fffffffffffff50003eb3c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf691c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ebc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b631c",
    x"070a0000000000000155fffffffffffff9ef35ea9a1c",
    x"08020000000000000155fffffffffffff6f669d9821c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2391c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee1a1c",
    x"0209000000000000015500000000000000fb335c1e1c",
    x"030b0000000000000155fffffffffffff50003eb3c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf661c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2eb81c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b5d1c",
    x"070a0000000000000155fffffffffffff9ef35ea961c",
    x"08020000000000000155fffffffffffff6f669d9801c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2351c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee1b1c",
    x"0209000000000000015500000000000000fb335c181c",
    x"030b0000000000000155fffffffffffff50003eb3d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf641c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2eb41c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b561c",
    x"070a0000000000000155fffffffffffff9ef35ea921c",
    x"08020000000000000155fffffffffffff6f669d97d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2311c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee1d1c",
    x"0209000000000000015500000000000000fb335c131c",
    x"030b0000000000000155fffffffffffff50003eb3e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf611c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2eb11c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b501c",
    x"070a0000000000000155fffffffffffff9ef35ea8e1c",
    x"08020000000000000155fffffffffffff6f669d97b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c22d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee1e1c",
    x"0209000000000000015500000000000000fb335c0d1c",
    x"030b0000000000000155fffffffffffff50003eb3f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf5e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2ead1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b4a1c",
    x"070a0000000000000155fffffffffffff9ef35ea8b1c",
    x"08020000000000000155fffffffffffff6f669d9781c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2291c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee1f1c",
    x"0209000000000000015500000000000000fb335c071c",
    x"030b0000000000000155fffffffffffff50003eb401c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf5c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2eaa1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b441c",
    x"070a0000000000000155fffffffffffff9ef35ea871c",
    x"08020000000000000155fffffffffffff6f669d9761c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c2241c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbee201c",
    x"0209000000000000031f00000000000000fb335c021c",
    x"030b000000000000031ffffffffffffff50003eb411c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbf591c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2ea61c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0b3e1c",
    x"070a000000000000031ffffffffffffff9ef35ea831c",
    x"0802000000000000031ffffffffffffff6f669d9741c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c2201c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbee211c",
    x"020900000000000000ae00000000000000fb335bfc1c",
    x"030b00000000000000aefffffffffffff50003eb421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbf571c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2ea31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0b381c",
    x"070a00000000000000aefffffffffffff9ef35ea7f1c",
    x"080200000000000000aefffffffffffff6f669d9711c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c21c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbee221c",
    x"020900000000000001a400000000000000fb335bf71c",
    x"030b00000000000001a4fffffffffffff50003eb421c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbf541c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2e9f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0b311c",
    x"070a00000000000001a4fffffffffffff9ef35ea7c1c",
    x"080200000000000001a4fffffffffffff6f669d96f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a6ffffffffffffff0266c2181c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a60000000000000b0bfbee231c",
    x"020900000000000001a600000000000000fb335bf11c",
    x"030b00000000000001a6fffffffffffff50003eb431c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a6fffffffffffff4099dbf521c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a60000000000000b072f2e9b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a60000000000000004cd0b2b1c",
    x"070a00000000000001a6fffffffffffff9ef35ea781c",
    x"080200000000000001a6fffffffffffff6f669d96c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2141c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee251c",
    x"0209000000000000015500000000000000fb335beb1c",
    x"030b0000000000000155fffffffffffff50003eb441c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf4f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e981c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b251c",
    x"070a0000000000000155fffffffffffff9ef35ea741c",
    x"08020000000000000155fffffffffffff6f669d96a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2101c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee261c",
    x"0209000000000000015500000000000000fb335be61c",
    x"030b0000000000000155fffffffffffff50003eb451c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf4d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e941c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b1f1c",
    x"070a0000000000000155fffffffffffff9ef35ea701c",
    x"08020000000000000155fffffffffffff6f669d9671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c20c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee271c",
    x"0209000000000000015500000000000000fb335be01c",
    x"030b0000000000000155fffffffffffff50003eb461c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf4a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e911c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b191c",
    x"070a0000000000000155fffffffffffff9ef35ea6d1c",
    x"08020000000000000155fffffffffffff6f669d9651c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2071c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee281c",
    x"0209000000000000015500000000000000fb335bdb1c",
    x"030b0000000000000155fffffffffffff50003eb471c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf471c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e8d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b121c",
    x"070a0000000000000155fffffffffffff9ef35ea691c",
    x"08020000000000000155fffffffffffff6f669d9631c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c2031c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee291c",
    x"0209000000000000015500000000000000fb335bd51c",
    x"030b0000000000000155fffffffffffff50003eb481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf451c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e891c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b0c1c",
    x"070a0000000000000155fffffffffffff9ef35ea651c",
    x"08020000000000000155fffffffffffff6f669d9601c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1ff1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee2a1c",
    x"0209000000000000015500000000000000fb335bcf1c",
    x"030b0000000000000155fffffffffffff50003eb481c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf421c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e861c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b061c",
    x"070a0000000000000155fffffffffffff9ef35ea611c",
    x"08020000000000000155fffffffffffff6f669d95e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1fb1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee2c1c",
    x"0209000000000000015500000000000000fb335bca1c",
    x"030b0000000000000155fffffffffffff50003eb491c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf401c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e821c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0b001c",
    x"070a0000000000000155fffffffffffff9ef35ea5e1c",
    x"08020000000000000155fffffffffffff6f669d95b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1f71c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee2d1c",
    x"0209000000000000015500000000000000fb335bc41c",
    x"030b0000000000000155fffffffffffff50003eb4a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf3d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e7f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0afa1c",
    x"070a0000000000000155fffffffffffff9ef35ea5a1c",
    x"08020000000000000155fffffffffffff6f669d9591c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1f31c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee2e1c",
    x"0209000000000000015500000000000000fb335bbe1c",
    x"030b0000000000000155fffffffffffff50003eb4b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf3b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e7b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0af31c",
    x"070a0000000000000155fffffffffffff9ef35ea561c",
    x"08020000000000000155fffffffffffff6f669d9561c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1ee1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee2f1c",
    x"0209000000000000015500000000000000fb335bb91c",
    x"030b0000000000000155fffffffffffff50003eb4c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf381c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e781c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0aed1c",
    x"070a0000000000000155fffffffffffff9ef35ea521c",
    x"08020000000000000155fffffffffffff6f669d9541c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1ea1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee301c",
    x"0209000000000000015500000000000000fb335bb31c",
    x"030b0000000000000155fffffffffffff50003eb4d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf361c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e741c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ae71c",
    x"070a0000000000000155fffffffffffff9ef35ea4f1c",
    x"08020000000000000155fffffffffffff6f669d9521c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1e61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee311c",
    x"0209000000000000015500000000000000fb335bae1c",
    x"030b0000000000000155fffffffffffff50003eb4e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf331c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e701c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ae11c",
    x"070a0000000000000155fffffffffffff9ef35ea4b1c",
    x"08020000000000000155fffffffffffff6f669d94f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1e21c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee321c",
    x"0209000000000000015500000000000000fb335ba81c",
    x"030b0000000000000155fffffffffffff50003eb4e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf311c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e6d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0adb1c",
    x"070a0000000000000155fffffffffffff9ef35ea471c",
    x"08020000000000000155fffffffffffff6f669d94d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1de1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee341c",
    x"0209000000000000015500000000000000fb335ba21c",
    x"030b0000000000000155fffffffffffff50003eb4f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf2e1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e691c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0ad41c",
    x"070a0000000000000155fffffffffffff9ef35ea431c",
    x"08020000000000000155fffffffffffff6f669d94a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c1da1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbee351c",
    x"0209000000000000029500000000000000fb335b9d1c",
    x"030b0000000000000295fffffffffffff50003eb501c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dbf2b1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f2e661c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd0ace1c",
    x"070a0000000000000295fffffffffffff9ef35ea401c",
    x"08020000000000000295fffffffffffff6f669d9481c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1d61c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee361c",
    x"020900000000000002aa00000000000000fb335b971c",
    x"030b00000000000002aafffffffffffff50003eb511c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbf291c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2e621c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0ac81c",
    x"070a00000000000002aafffffffffffff9ef35ea3c1c",
    x"080200000000000002aafffffffffffff6f669d9451c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c1d11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbee371c",
    x"0209000000000000031f00000000000000fb335b911c",
    x"030b000000000000031ffffffffffffff50003eb521c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbf261c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2e5f1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0ac21c",
    x"070a000000000000031ffffffffffffff9ef35ea381c",
    x"0802000000000000031ffffffffffffff6f669d9431c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c1cd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbee381c",
    x"020900000000000000ae00000000000000fb335b8c1c",
    x"030b00000000000000aefffffffffffff50003eb531c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbf241c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2e5b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0abc1c",
    x"070a00000000000000aefffffffffffff9ef35ea341c",
    x"080200000000000000aefffffffffffff6f669d9411c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c1c91c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbee391c",
    x"020900000000000001a400000000000000fb335b861c",
    x"030b00000000000001a4fffffffffffff50003eb541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbf211c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2e571c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0ab51c",
    x"070a00000000000001a4fffffffffffff9ef35ea311c",
    x"080200000000000001a4fffffffffffff6f669d93e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000166ffffffffffffff0266c1c51c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001660000000000000b0bfbee3a1c",
    x"0209000000000000016600000000000000fb335b811c",
    x"030b0000000000000166fffffffffffff50003eb541c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000166fffffffffffff4099dbf1f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001660000000000000b072f2e541c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001660000000000000004cd0aaf1c",
    x"070a0000000000000166fffffffffffff9ef35ea2d1c",
    x"08020000000000000166fffffffffffff6f669d93c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000295ffffffffffffff0266c1c11c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002950000000000000b0bfbee3c1c",
    x"0209000000000000029500000000000000fb335b7b1c",
    x"030b0000000000000295fffffffffffff50003eb551c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000295fffffffffffff4099dbf1c1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002950000000000000b072f2e501c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002950000000000000004cd0aa91c",
    x"070a0000000000000295fffffffffffff9ef35ea291c",
    x"08020000000000000295fffffffffffff6f669d9391c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000159ffffffffffffff0266c1bd1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001590000000000000b0bfbee3d1c",
    x"0209000000000000015900000000000000fb335b751c",
    x"030b0000000000000159fffffffffffff50003eb561c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000159fffffffffffff4099dbf1a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001590000000000000b072f2e4d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001590000000000000004cd0aa31c",
    x"070a0000000000000159fffffffffffff9ef35ea251c",
    x"08020000000000000159fffffffffffff6f669d9371c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1b81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee3e1c",
    x"0209000000000000015500000000000000fb335b701c",
    x"030b0000000000000155fffffffffffff50003eb571c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf171c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e491c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a9d1c",
    x"070a0000000000000155fffffffffffff9ef35ea221c",
    x"08020000000000000155fffffffffffff6f669d9341c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1b41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee3f1c",
    x"0209000000000000015500000000000000fb335b6a1c",
    x"030b0000000000000155fffffffffffff50003eb581c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf141c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e461c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a961c",
    x"070a0000000000000155fffffffffffff9ef35ea1e1c",
    x"08020000000000000155fffffffffffff6f669d9321c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1b01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee401c",
    x"0209000000000000015500000000000000fb335b641c",
    x"030b0000000000000155fffffffffffff50003eb591c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf121c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e421c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a901c",
    x"070a0000000000000155fffffffffffff9ef35ea1a1c",
    x"08020000000000000155fffffffffffff6f669d9301c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1ac1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee411c",
    x"0209000000000000015500000000000000fb335b5f1c",
    x"030b0000000000000155fffffffffffff50003eb5a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf0f1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e3e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a8a1c",
    x"070a0000000000000155fffffffffffff9ef35ea161c",
    x"08020000000000000155fffffffffffff6f669d92d1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1a81c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee421c",
    x"0209000000000000015500000000000000fb335b591c",
    x"030b0000000000000155fffffffffffff50003eb5a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf0d1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e3b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a841c",
    x"070a0000000000000155fffffffffffff9ef35ea121c",
    x"08020000000000000155fffffffffffff6f669d92b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1a41c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee441c",
    x"0209000000000000015500000000000000fb335b541c",
    x"030b0000000000000155fffffffffffff50003eb5b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf0a1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e371c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a7e1c",
    x"070a0000000000000155fffffffffffff9ef35ea0f1c",
    x"08020000000000000155fffffffffffff6f669d9281c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1a01c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee451c",
    x"0209000000000000015500000000000000fb335b4e1c",
    x"030b0000000000000155fffffffffffff50003eb5c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf081c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e341c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a771c",
    x"070a0000000000000155fffffffffffff9ef35ea0b1c",
    x"08020000000000000155fffffffffffff6f669d9261c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c19b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee461c",
    x"0209000000000000015500000000000000fb335b481c",
    x"030b0000000000000155fffffffffffff50003eb5d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf051c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e301c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a711c",
    x"070a0000000000000155fffffffffffff9ef35ea071c",
    x"08020000000000000155fffffffffffff6f669d9231c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1971c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee471c",
    x"0209000000000000015500000000000000fb335b431c",
    x"030b0000000000000155fffffffffffff50003eb5e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf031c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e2d1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a6b1c",
    x"070a0000000000000155fffffffffffff9ef35ea031c",
    x"08020000000000000155fffffffffffff6f669d9211c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1931c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee481c",
    x"0209000000000000015500000000000000fb335b3d1c",
    x"030b0000000000000155fffffffffffff50003eb5f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbf001c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e291c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a651c",
    x"070a0000000000000155fffffffffffff9ef35ea001c",
    x"08020000000000000155fffffffffffff6f669d91f1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c18f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee491c",
    x"0209000000000000015500000000000000fb335b371c",
    x"030b0000000000000155fffffffffffff50003eb5f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbefd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e251c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a5f1c",
    x"070a0000000000000155fffffffffffff9ef35e9fc1c",
    x"08020000000000000155fffffffffffff6f669d91c1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c18b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee4b1c",
    x"0209000000000000015500000000000000fb335b321c",
    x"030b0000000000000155fffffffffffff50003eb601c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbefb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e221c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a581c",
    x"070a0000000000000155fffffffffffff9ef35e9f81c",
    x"08020000000000000155fffffffffffff6f669d91a1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000255ffffffffffffff0266c1871c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002550000000000000b0bfbee4c1c",
    x"0209000000000000025500000000000000fb335b2c1c",
    x"030b0000000000000255fffffffffffff50003eb611c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000255fffffffffffff4099dbef81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002550000000000000b072f2e1e1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002550000000000000004cd0a521c",
    x"070a0000000000000255fffffffffffff9ef35e9f41c",
    x"08020000000000000255fffffffffffff6f669d9171c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000155ffffffffffffff0266c1831c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001550000000000000b0bfbee4d1c",
    x"0209000000000000015500000000000000fb335b271c",
    x"030b0000000000000155fffffffffffff50003eb621c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000155fffffffffffff4099dbef61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001550000000000000b072f2e1b1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001550000000000000004cd0a4c1c",
    x"070a0000000000000155fffffffffffff9ef35e9f11c",
    x"08020000000000000155fffffffffffff6f669d9151c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c17e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbee4e1c",
    x"0209000000000000031f00000000000000fb335b211c",
    x"030b000000000000031ffffffffffffff50003eb631c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbef31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2e171c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd0a461c",
    x"070a000000000000031ffffffffffffff9ef35e9ed1c",
    x"0802000000000000031ffffffffffffff6f669d9121c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c17a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbee4f1c",
    x"020900000000000000ae00000000000000fb335b1b1c",
    x"030b00000000000000aefffffffffffff50003eb641c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbef11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2e141c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd0a401c",
    x"070a00000000000000aefffffffffffff9ef35e9e91c",
    x"080200000000000000aefffffffffffff6f669d9101c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c1761c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbee501c",
    x"020900000000000001a400000000000000fb335b161c",
    x"030b00000000000001a4fffffffffffff50003eb651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbeee1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2e101c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd0a3a1c",
    x"070a00000000000001a4fffffffffffff9ef35e9e51c",
    x"080200000000000001a4fffffffffffff6f669d90e1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"00010000000000000266ffffffffffffff0266c1721c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002660000000000000b0bfbee511c",
    x"0209000000000000026600000000000000fb335b101c",
    x"030b0000000000000266fffffffffffff50003eb651c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"04110000000000000266fffffffffffff4099dbeec1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002660000000000000b072f2e0c1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002660000000000000004cd0a331c",
    x"070a0000000000000266fffffffffffff9ef35e9e21c",
    x"08020000000000000266fffffffffffff6f669d90b1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c16e1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee531c",
    x"020900000000000002aa00000000000000fb335b0a1c",
    x"030b00000000000002aafffffffffffff50003eb661c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbee91c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2e091c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a2d1c",
    x"070a00000000000002aafffffffffffff9ef35e9de1c",
    x"080200000000000002aafffffffffffff6f669d9091c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c16a1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee541c",
    x"020900000000000002aa00000000000000fb335b051c",
    x"030b00000000000002aafffffffffffff50003eb671c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbee61c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2e051c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a271c",
    x"070a00000000000002aafffffffffffff9ef35e9da1c",
    x"080200000000000002aafffffffffffff6f669d9061c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1651c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee551c",
    x"020900000000000002aa00000000000000fb335aff1c",
    x"030b00000000000002aafffffffffffff50003eb681c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbee41c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2e021c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a211c",
    x"070a00000000000002aafffffffffffff9ef35e9d61c",
    x"080200000000000002aafffffffffffff6f669d9041c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1611c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee561c",
    x"020900000000000002aa00000000000000fb335afa1c",
    x"030b00000000000002aafffffffffffff50003eb691c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbee11c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dfe1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a1b1c",
    x"070a00000000000002aafffffffffffff9ef35e9d31c",
    x"080200000000000002aafffffffffffff6f669d9011c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c15d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee571c",
    x"020900000000000002aa00000000000000fb335af41c",
    x"030b00000000000002aafffffffffffff50003eb6a1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbedf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dfb1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a141c",
    x"070a00000000000002aafffffffffffff9ef35e9cf1c",
    x"080200000000000002aafffffffffffff6f669d8ff1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1591c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee581c",
    x"020900000000000002aa00000000000000fb335aee1c",
    x"030b00000000000002aafffffffffffff50003eb6b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbedc1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2df71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a0e1c",
    x"070a00000000000002aafffffffffffff9ef35e9cb1c",
    x"080200000000000002aafffffffffffff6f669d8fd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1551c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee591c",
    x"020900000000000002aa00000000000000fb335ae91c",
    x"030b00000000000002aafffffffffffff50003eb6b1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbeda1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2df31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a081c",
    x"070a00000000000002aafffffffffffff9ef35e9c71c",
    x"080200000000000002aafffffffffffff6f669d8fa1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1511c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee5b1c",
    x"020900000000000002aa00000000000000fb335ae31c",
    x"030b00000000000002aafffffffffffff50003eb6c1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbed71c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2df01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd0a021c",
    x"070a00000000000002aafffffffffffff9ef35e9c41c",
    x"080200000000000002aafffffffffffff6f669d8f81c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c14d1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee5c1c",
    x"020900000000000002aa00000000000000fb335add1c",
    x"030b00000000000002aafffffffffffff50003eb6d1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbed51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dec1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09fc1c",
    x"070a00000000000002aafffffffffffff9ef35e9c01c",
    x"080200000000000002aafffffffffffff6f669d8f51c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1481c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee5d1c",
    x"020900000000000002aa00000000000000fb335ad81c",
    x"030b00000000000002aafffffffffffff50003eb6e1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbed21c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2de91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09f51c",
    x"070a00000000000002aafffffffffffff9ef35e9bc1c",
    x"080200000000000002aafffffffffffff6f669d8f31c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1441c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee5e1c",
    x"020900000000000002aa00000000000000fb335ad21c",
    x"030b00000000000002aafffffffffffff50003eb6f1c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbecf1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2de51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09ef1c",
    x"070a00000000000002aafffffffffffff9ef35e9b81c",
    x"080200000000000002aafffffffffffff6f669d8f01c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1401c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee5f1c",
    x"020900000000000002aa00000000000000fb335acd1c",
    x"030b00000000000002aafffffffffffff50003eb701c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbecd1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2de21c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09e91c",
    x"070a00000000000002aafffffffffffff9ef35e9b41c",
    x"080200000000000002aafffffffffffff6f669d8ee1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c13c1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee601c",
    x"020900000000000002aa00000000000000fb335ac71c",
    x"030b00000000000002aafffffffffffff50003eb711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbeca1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dde1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09e31c",
    x"070a00000000000002aafffffffffffff9ef35e9b11c",
    x"080200000000000002aafffffffffffff6f669d8ec1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1381c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee621c",
    x"020900000000000002aa00000000000000fb335ac11c",
    x"030b00000000000002aafffffffffffff50003eb711c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbec81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dda1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09dd1c",
    x"070a00000000000002aafffffffffffff9ef35e9ad1c",
    x"080200000000000002aafffffffffffff6f669d8e91c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1341c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee631c",
    x"020900000000000002aa00000000000000fb335abc1c",
    x"030b00000000000002aafffffffffffff50003eb721c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbec51c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dd71c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09d61c",
    x"070a00000000000002aafffffffffffff9ef35e9a91c",
    x"080200000000000002aafffffffffffff6f669d8e71c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000002aaffffffffffffff0266c1301c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000002aa0000000000000b0bfbee641c",
    x"020900000000000002aa00000000000000fb335ab61c",
    x"030b00000000000002aafffffffffffff50003eb731c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000002aafffffffffffff4099dbec31c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000002aa0000000000000b072f2dd31c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000002aa0000000000000004cd09d01c",
    x"070a00000000000002aafffffffffffff9ef35e9a51c",
    x"080200000000000002aafffffffffffff6f669d8e41c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"0001000000000000031fffffffffffffff0266c12b1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"0107000000000000031f0000000000000b0bfbee651c",
    x"0209000000000000031f00000000000000fb335ab01c",
    x"030b000000000000031ffffffffffffff50003eb741c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"0411000000000000031ffffffffffffff4099dbec01c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"0517000000000000031f0000000000000b072f2dd01c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"0618000000000000031f0000000000000004cd09ca1c",
    x"070a000000000000031ffffffffffffff9ef35e9a21c",
    x"0802000000000000031ffffffffffffff6f669d8e21c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000000aeffffffffffffff0266c1271c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000000ae0000000000000b0bfbee661c",
    x"020900000000000000ae00000000000000fb335aab1c",
    x"030b00000000000000aefffffffffffff50003eb751c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000000aefffffffffffff4099dbebe1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000000ae0000000000000b072f2dcc1c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000000ae0000000000000004cd09c41c",
    x"070a00000000000000aefffffffffffff9ef35e99e1c",
    x"080200000000000000aefffffffffffff6f669d8df1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001a4ffffffffffffff0266c1231c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001a40000000000000b0bfbee671c",
    x"020900000000000001a400000000000000fb335aa51c",
    x"030b00000000000001a4fffffffffffff50003eb761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001a4fffffffffffff4099dbebb1c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001a40000000000000b072f2dc91c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001a40000000000000004cd09be1c",
    x"070a00000000000001a4fffffffffffff9ef35e99a1c",
    x"080200000000000001a4fffffffffffff6f669d8dd1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"000100000000000001aaffffffffffffff0266c11f1c",
    x"ffff0000000000000000000000000000000c0000001c",
    x"ffff000000000000000000000000000000026666661c",
    x"010700000000000001aa0000000000000b0bfbee681c",
    x"020900000000000001aa00000000000000fb335aa01c",
    x"030b00000000000001aafffffffffffff50003eb761c",
    x"ffff000000000000000000000000000000fb3333341c",
    x"ffff000000000000000000000000000000000000001c",
    x"041100000000000001aafffffffffffff4099dbeb81c",
    x"ffff000000000000000000000000000000073333331c",
    x"ffff000000000000000000000000000000099999991c",
    x"051700000000000001aa0000000000000b072f2dc51c",
    x"ffff000000000000000000000000000000f66666671c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"061800000000000001aa0000000000000004cd09b71c",
    x"070a00000000000001aafffffffffffff9ef35e9961c",
    x"080200000000000001aafffffffffffff6f669d8da1c",
    x"ffff000000000000000000000000000000fd99999a1c",
    x"ffff000000000000000000000000000000f8cccccd1c",
    x"ffff0000000000000000000000000000000e6666661c",
    x"ffff000000000000000000000000000000ef3333341c",
    x"ffff00000000000000000000000000000004cccccc1c",
    x"ffff000000000000000000000000000000f8cccccd1c"
  );
end package;