library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package input is
  
  constant inputFrameSatCount : integer := 1;
  
  type inputTable is array(0 to 100 - 1) of std_logic_vector(176-1 downto 0);
  constant inputSeq : inputTable := (
    x"000100000000000000110000000271411afffeee76ff",
    x"00010000000000000006ffffffffffffe5fffeee63ff",
    x"000100000000000000000000000000000afffeee4fff",
    x"000100000000000000000000000000000bfffeee3cff",
    x"000100000000000000140000000000000bfffeee28ff",
    x"0001000000000000001d0000000000000bfffeee15ff",
    x"000100000000000000050000000000000bfffeee01ff",
    x"0001000000000000001b0000000000000bfffeedeeff",
    x"0001000000000000001d0000000000000cfffeeddaff",
    x"0001000000000000001d0000000000000bfffeedc7ff",
    x"0001000000000000001d0000000000000bfffeedb3ff",
    x"000100000000000000000000000000000bfffeeda0ff",
    x"0001000000000000001c0000000000000bfffeed8cff",
    x"000100000000000000110000000000000bfffeed79ff",
    x"000100000000000000020000000000000bfffeed65ff",
    x"0001000000000000001e0000000000000bfffeed52ff",
    x"000100000000000000030000000000000bfffeed3eff",
    x"000100000000000000030000000000000bfffeed2bff",
    x"000100000000000000000000000000000bfffeed17ff",
    x"000100000000000000000000000000000bfffeed04ff",
    x"000100000000000000000000000000000bfffeecf0ff",
    x"000100000000000000000000000000000bfffeecddff",
    x"000100000000000000000000000000000bfffeecc9ff",
    x"000100000000000000000000000000000bfffeecb6ff",
    x"000100000000000000000000000000000cfffeeca2ff",
    x"000100000000000000000000000000000bfffeec8fff",
    x"000100000000000000000000000000000bfffeec7bff",
    x"000100000000000000000000000000000bfffeec68ff",
    x"000100000000000000000000000000000bfffeec54ff",
    x"000100000000000000000000000000000bfffeec41ff",
    x"000100000000000000000000000000000bfffeec2dff",
    x"000100000000000000000000000000000bfffeec1aff",
    x"000100000000000000000000000000000bfffeec06ff",
    x"000100000000000000000000000000000bfffeebf3ff",
    x"000100000000000000000000000000000cfffeebdfff",
    x"000100000000000000000000000000000bfffeebccff",
    x"000100000000000000000000000000000bfffeebb8ff",
    x"000100000000000000000000000000000bfffeeba5ff",
    x"000100000000000000000000000000000bfffeeb91ff",
    x"000100000000000000000000000000000bfffeeb7dff",
    x"0001000000000000001d0000000000000bfffeeb6aff",
    x"000100000000000000000000000000000bfffeeb57ff",
    x"0001000000000000001a0000000000000cfffeeb43ff",
    x"000100000000000000020000000000000bfffeeb2fff",
    x"000100000000000000000000000000000bfffeeb1cff",
    x"000100000000000000000000000000000bfffeeb08ff",
    x"000100000000000000000000000000000bfffeeaf5ff",
    x"000100000000000000170000000000000bfffeeae1ff",
    x"0001000000000000001f0000000000000bfffeeaceff",
    x"0001000000000000001f0000000000000cfffeeabaff",
    x"0001000000000000001f0000000000000bfffeeaa7ff",
    x"0001000000000000001f0000000000000bfffeea93ff",
    x"0001000000000000001b0000000000000bfffeea80ff",
    x"000100000000000000190000000000000bfffeea6cff",
    x"000100000000000000170000000000000cfffeea59ff",
    x"0001000000000000000a0000000000000bfffeea45ff",
    x"000100000000000000060000000000000bfffeea32ff",
    x"0001000000000000000f0000000000000bfffeea1eff",
    x"000100000000000000040000000000000bfffeea0bff",
    x"000100000000000000020000000000000bfffee9f7ff",
    x"000100000000000000110000000000000cfffee9e4ff",
    x"000100000000000000060000000000000bfffee9d0ff",
    x"000100000000000000000000000000000bfffee9bdff",
    x"000100000000000000000000000000000bfffee9a9ff",
    x"000100000000000000140000000000000bfffee996ff",
    x"0001000000000000001d0000000000000cfffee982ff",
    x"000100000000000000050000000000000bfffee96fff",
    x"0001000000000000001b0000000000000bfffee95bff",
    x"0001000000000000001d0000000000000bfffee948ff",
    x"0001000000000000001e0000000000000cfffee934ff",
    x"0001000000000000001a0000000000000bfffee921ff",
    x"000100000000000000010000000000000bfffee90dff",
    x"0001000000000000001a0000000000000bfffee8faff",
    x"000100000000000000020000000000000bfffee8e6ff",
    x"000100000000000000000000000000000cfffee8d3ff",
    x"0001000000000000000d0000000000000bfffee8bfff",
    x"000100000000000000070000000000000bfffee8acff",
    x"000100000000000000000000000000000bfffee898ff",
    x"000100000000000000140000000000000cfffee885ff",
    x"000100000000000000120000000000000bfffee871ff",
    x"000100000000000000120000000000000bfffee85eff",
    x"000100000000000000090000000000000bfffee84aff",
    x"0001000000000000001e0000000000000cfffee836ff",
    x"000100000000000000000000000000000bfffee823ff",
    x"0001000000000000001d0000000000000bfffee80fff",
    x"0001000000000000001f0000000000000cfffee7fcff",
    x"000100000000000000070000000000000bfffee7e8ff",
    x"000100000000000000080000000000000bfffee7d5ff",
    x"0001000000000000001f0000000000000bfffee7c1ff",
    x"000100000000000000000000000000000cfffee7aeff",
    x"000100000000000000000000000000000bfffee79aff",
    x"000100000000000000140000000000000bfffee787ff",
    x"0001000000000000001b0000000000000cfffee773ff",
    x"000100000000000000010000000000000bfffee760ff",
    x"000100000000000000160000000000000bfffee74cff",
    x"0001000000000000000c0000000000000bfffee739ff",
    x"000100000000000000050000000000000cfffee725ff",
    x"000100000000000000060000000000000bfffee712ff",
    x"0001000000000000001c0000000000000bfffee6feff",
    x"000100000000000000040000000000000cfffee6ebff"
  );
end package;