library ieee;
use ieee.std_logic_1164.all;
USE ieee.std_logic_arith.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
library std;
use STD.textio.all;
use work.settings.all;


entity InputHandler_tb is
end;

architecture bench of InputHandler_tb is
    
    --constant frameWidth: integer := 176;
    --constant chanel_count : integer := 4;

    component SPI_helper
        generic (
          n : integer := frameWidth;
          clk_period : time := samplePeriode
        );
        port (
          word : in std_logic_vector(frameWidth-1 downto 0);
          done : out std_logic;
          clk : out std_logic;
          serial_out : out std_logic
        );
    end component;
    
    component InputHandler
        generic (
          chanel_count : integer := chanel_count
        );
        port (
          clk : in std_logic;
          reset : in std_logic;
          serial_in : in std_logic;
          store : in std_logic;
          I : out IQ;
          Q : out IQ
        );
    end component;

    signal clk       : std_logic := '0';
    signal reset     : std_logic := '0';
    signal send_done : std_logic := '0';
    signal serial    : std_logic := '0';
    signal store     : std_logic := '0';

    signal I, Q : IQ;

    signal word    : std_logic_vector(frameWidth-1 downto 0);

    file IQ_file : text;
    signal sim_running : boolean := false;
    signal sim_stopping : boolean := false;
begin

    InputHandler0: InputHandler port map (clk, reset, serial, store, I, Q);
    SPI_HELPER0: SPI_helper port map (word, send_done, clk, serial);

    reset <= '1', '0' after 1 ns;

    process
    begin
      wait for 15000 ms;
      sim_stopping <= true;
    end process;


    process
      variable iqLine     : line;
    begin
      wait for 90 ms;
      sim_running <= true;
      wait for 1 ms;
      file_open(IQ_file, "output_results.txt", write_mode);
      while sim_running=true or sim_stopping=false loop
        wait until falling_edge(clk);
        write(iqLine, to_integer(I));
        write(iqLine, string'(", "));
        write(iqLine, to_integer(Q));
        writeline(IQ_file, iqLine);
        wait for 25 ns;
      end loop;
    file_close(IQ_file);
    report "done";
    wait;
    end process;

    process

        procedure send(value: in std_logic_vector(frameWidth-1 downto 0)) is
        begin
            word <= value;
            wait until rising_edge(send_done);
            store <= '1';
            wait for 0.5 us;
            store <= '0';
            wait for 0.5 us;
        end procedure;

        procedure send(
          satNum:     in integer range 0 to 255;
          bits:       in std_logic_vector(63 downto 0);
          delay:      in std_logic_vector(63 downto 0);
          phase_step: in integer;
          power:      in integer range 0 to 255
        ) is
        begin
            send(
              std_logic_vector(to_unsigned(satNum, 8)) & 
              bits & 
              delay & 
              std_logic_vector(to_signed(phase_step, 32)) & 
              std_logic_vector(to_unsigned(power, 8))
            );
        end procedure;

        procedure send(
          satNum:     in integer range 0 to 255;
          bits:       in std_logic_vector(63 downto 0);
          delay:      in integer;
          phase_step: in integer;
          power:      in integer range 0 to 255
        ) is
        begin
            send(
              satNum, bits,
              std_logic_vector(to_signed(delay, 64)),
              phase_step, power
            );
        end procedure;

    begin
        wait for 1 us;
        --send(x"00333333333333333333333333333333333333333333");
        --send(0, x"3333333333333333", 0, 10, 255);
        --wait for 10 us;
        --send(x"01aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa");
        --send(1, x"aaaaaaaaaaaaaaaa", 0, 20, 0);
        --wait for 10 us;
        --send(x"02555555555555555555555555555555555555555555");
        --send(2, x"5555555555555555", 0, 0, 0);
        --wait for 10 us;
        --send(x"03999999999999999999999999999999999999999999");
        --send(3, x"9999999999999999", 0, 0, 0);
        --wait for 10 us;

        send(0, x"00000000000001aa", x"00002d0fe08c7ccf", 40297315, 62);
send(1, x"00000000000001aa", x"0000376488083bd7", -80508804, 62);
send(2, x"00000000000001aa", x"000033b172389eb7", 161338012, 62);
send(3, x"00000000000001aa", x"000030e7165c8831", 120540046, 62);
send(0, x"0000000000000295", x"00002d0fdf463844", 40297315, 62);
send(1, x"0000000000000295", x"000037648729259a", -80508804, 62);
send(2, x"0000000000000295", x"000033b167359ff8", 161338012, 62);
send(3, x"0000000000000295", x"000030e7208b4546", 120540046, 62);
send(0, x"000000000000015a", x"00002d0fddffffb2", 40297244, 62);
send(1, x"000000000000015a", x"00003764864a1858", -80508804, 62);
send(2, x"000000000000015a", x"000033b15c32a13a", 161338012, 62);
send(3, x"000000000000015a", x"000030e72aba0e54", 120540046, 62);
send(0, x"0000000000000155", x"00002d0fdcb9d01b", 40297244, 62);
send(1, x"0000000000000155", x"00003764856b1d0e", -80508804, 62);
send(2, x"0000000000000155", x"000033b1512fae76", 161338012, 62);
send(3, x"0000000000000155", x"000030e734e8e05f", 120540046, 62);
send(0, x"00000000000001a9", x"00002d0fdb73af7d", 40297244, 62);
send(1, x"00000000000002a9", x"00003764848c2dbd", -80508804, 62);
send(2, x"0000000000000295", x"000033b1462cc1ae", 161338012, 62);
send(3, x"0000000000000155", x"000030e73f17bb64", 120540046, 62);
send(0, x"00000000000002a6", x"00002d0fda2d94dc", 40297244, 62);
send(1, x"000000000000029a", x"0000376483ad5064", -80508804, 62);
send(2, x"0000000000000165", x"000033b13b29d7e5", 161338012, 62);
send(3, x"0000000000000256", x"000030e74946a264", 120540046, 62);
send(0, x"000000000000016a", x"00002d0fd8e78635", 40297244, 62);
send(1, x"000000000000015a", x"0000376482ce7f04", -80508875, 62);
send(2, x"0000000000000196", x"000033b13026f419", 161338012, 62);
send(3, x"00000000000002aa", x"000030e75375925f", 120540046, 62);
send(0, x"00000000000001a9", x"00002d0fd7a18388", 40297244, 62);
send(1, x"0000000000000199", x"0000376481efbc9d", -80508875, 62);
send(2, x"000000000000025a", x"000033b125241948", 161338012, 62);
send(3, x"00000000000001a6", x"000030e75da48b55", 120540046, 62);
send(0, x"0000000000000266", x"00002d0fd65b8cd5", 40297244, 62);
send(1, x"0000000000000166", x"000037648111092f", -80508875, 62);
send(2, x"0000000000000196", x"000033b11a214475", 161338012, 62);
send(3, x"0000000000000259", x"000030e767d38d47", 120540046, 62);
send(0, x"000000000000025a", x"00002d0fd515a21c", 40297244, 62);
send(1, x"0000000000000155", x"00003764803264b9", -80508875, 62);
send(2, x"00000000000001a5", x"000033b10f1e72a0", 161338012, 62);
send(3, x"000000000000016a", x"000030e772029b33", 120540046, 62);
send(0, x"0000000000000256", x"00002d0fd3cfc05f", 40297244, 62);
send(1, x"000000000000015a", x"000037647f53cf3b", -80508875, 62);
send(2, x"00000000000002aa", x"000033b1041ba9c7", 161338012, 62);
send(3, x"0000000000000269", x"000030e77c31b21a", 120540046, 62);
send(0, x"00000000000001a6", x"00002d0fd289ea9b", 40297244, 62);
send(1, x"00000000000001a9", x"000037647e7545b8", -80508875, 62);
send(2, x"0000000000000255", x"000033b0f918e3ec", 161338012, 62);
send(3, x"0000000000000156", x"000030e78660d1fe", 120540046, 62);
send(0, x"0000000000000196", x"00002d0fd14420d2", 40297244, 62);
send(1, x"00000000000002aa", x"000037647d96cb2d", -80508875, 62);
send(2, x"000000000000025a", x"000033b0ee16270c", 161338012, 62);
send(3, x"0000000000000295", x"000030e7908ffadc", 120540046, 62);
send(0, x"0000000000000299", x"00002d0fcffe6004", 40297244, 62);
send(1, x"000000000000029a", x"000037647cb86299", -80508875, 62);
send(2, x"00000000000002a5", x"000033b0e313702a", 161338012, 62);
send(3, x"0000000000000295", x"000030e79abf2fb4", 120540046, 62);
send(0, x"0000000000000199", x"00002d0fceb8ab30", 40297244, 62);
send(1, x"00000000000002a6", x"000037647bda05fe", -80508875, 62);
send(2, x"0000000000000269", x"000033b0d810bf44", 161338012, 62);
send(3, x"0000000000000295", x"000030e7a4ee6a8a", 120540046, 62);
send(0, x"0000000000000166", x"00002d0fcd72ff57", 40297244, 62);
send(1, x"000000000000015a", x"000037647afbbb5c", -80508875, 62);
send(2, x"000000000000016a", x"000033b0cd0e145c", 161338012, 62);
send(3, x"0000000000000299", x"000030e7af1db458", 120539975, 62);
send(0, x"00000000000002a6", x"00002d0fcc2d5f79", 40297244, 62);
send(1, x"00000000000002a6", x"000037647a1d79b4", -80508875, 62);
send(2, x"000000000000015a", x"000033b0c20b6c72", 161338012, 62);
send(3, x"00000000000002aa", x"000030e7b94d0721", 120539975, 62);
send(0, x"000000000000031f", x"00002d0fcae7cb94", 40297244, 62);
send(1, x"000000000000031f", x"00003764793f4a04", -80508875, 62);
send(2, x"000000000000031f", x"000033b0b708cd83", 161338012, 62);
send(3, x"000000000000031f", x"000030e7c37c5fe8", 120539975, 62);
send(0, x"00000000000000ae", x"00002d0fc9a240ab", 40297244, 62);
send(1, x"00000000000000ae", x"000037647861294c", -80508875, 62);
send(2, x"00000000000000ae", x"000033b0ac063492", 161338012, 62);
send(3, x"00000000000000ae", x"000030e7cdabc4a9", 120539975, 62);
send(0, x"00000000000001a4", x"00002d0fc85cc1bc", 40297172, 62);
send(1, x"00000000000001a4", x"000037647783148d", -80508947, 62);
send(2, x"00000000000001a4", x"000033b0a1039e9f", 161338012, 62);
send(3, x"00000000000001a4", x"000030e7d7db3265", 120539975, 62);
send(0, x"000000000000016a", x"00002d0fc7174ec7", 40297172, 62);
send(1, x"000000000000016a", x"0000376476a511c7", -80508947, 62);
send(2, x"000000000000016a", x"000033b0960114a6", 161338012, 62);
send(3, x"000000000000016a", x"000030e7e20aac1b", 120539975, 62);
send(0, x"0000000000000155", x"00002d0fc5d1e7cc", 40297172, 62);
send(1, x"0000000000000155", x"0000376475c71df8", -80508947, 62);
send(2, x"0000000000000155", x"000033b08afe8dab", 161337941, 62);
send(3, x"0000000000000155", x"000030e7ec3a2bce", 120539975, 62);
send(0, x"0000000000000195", x"00002d0fc48c89cd", 40297172, 62);
send(1, x"0000000000000195", x"0000376474e93325", -80508947, 62);
send(2, x"0000000000000195", x"000033b07ffc09af", 161337941, 62);
send(3, x"0000000000000195", x"000030e7f669b77b", 120539975, 62);
send(0, x"00000000000002aa", x"00002d0fc34737c7", 40297172, 62);
send(1, x"00000000000002aa", x"00003764740b5d48", -80508947, 62);
send(2, x"00000000000002aa", x"000033b074f991ad", 161337941, 62);
send(3, x"00000000000002aa", x"000030e800994c23", 120539975, 62);
send(0, x"00000000000001aa", x"00002d0fc201f1bc", 40297172, 62);
send(1, x"0000000000000296", x"00003764732d9364", -80508947, 62);
send(2, x"00000000000001aa", x"000033b069f71ca9", 161337941, 62);
send(3, x"00000000000002aa", x"000030e80ac8ecc6", 120539975, 62);
send(0, x"00000000000001a5", x"00002d0fc0bcb4ac", 40297172, 62);
send(1, x"0000000000000265", x"00003764724fd879", -80508947, 62);
send(2, x"0000000000000299", x"000033b05ef4b0a1", 161337941, 62);
send(3, x"000000000000015a", x"000030e814f89663", 120539975, 62);
send(0, x"0000000000000259", x"00002d0fbf778097", 40297172, 62);
send(1, x"0000000000000296", x"0000376471722988", -80508947, 62);
send(2, x"000000000000019a", x"000033b053f24499", 161337941, 62);
send(3, x"0000000000000156", x"000030e81f2848fd", 120539975, 62);
send(0, x"0000000000000159", x"00002d0fbe32587c", 40297172, 62);
send(1, x"0000000000000169", x"0000376470948c8e", -80508947, 62);
send(2, x"0000000000000269", x"000033b048efe48c", 161337941, 62);
send(3, x"0000000000000295", x"000030e829580492", 120539975, 62);
send(0, x"000000000000016a", x"00002d0fbced3f5b", 40297172, 62);
send(1, x"00000000000002a5", x"000037646fb6fe8d", -80508947, 62);
send(2, x"00000000000001a5", x"000033b03ded877c", 161337941, 62);
send(3, x"00000000000002a6", x"000030e83387cc21", 120539975, 62);
send(0, x"000000000000026a", x"00002d0fbba82f34", 40297172, 62);
send(1, x"0000000000000255", x"000037646ed97987", -80508947, 62);
send(2, x"00000000000001aa", x"000033b032eb3069", 161337941, 62);
send(3, x"00000000000002a5", x"000030e83db799ad", 120539975, 62);
send(0, x"0000000000000295", x"00002d0fba632809", 40297172, 62);
send(1, x"000000000000029a", x"000037646dfc0976", -80508947, 62);
send(2, x"000000000000025a", x"000033b027e8df54", 161337941, 62);
send(3, x"000000000000015a", x"000030e847e77333", 120539975, 62);
send(0, x"00000000000002aa", x"00002d0fb91e2fd7", 40297172, 62);
send(1, x"00000000000001a6", x"000037646d1ea55f", -80508947, 62);
send(2, x"0000000000000159", x"000033b01ce6973a", 161337941, 62);
send(3, x"000000000000026a", x"000030e8521758b3", 120539975, 62);
send(0, x"00000000000002a5", x"00002d0fb7d93da1", 40297172, 62);
send(1, x"000000000000025a", x"000037646c414d43", -80509018, 62);
send(2, x"000000000000016a", x"000033b011e4521e", 161337941, 62);
send(3, x"0000000000000166", x"000030e85c474430", 120539975, 62);
send(0, x"0000000000000256", x"00002d0fb6945a64", 40297172, 62);
send(1, x"0000000000000296", x"000037646b64071e", -80509018, 62);
send(2, x"0000000000000165", x"000033b006e215ff", 161337941, 62);
send(3, x"000000000000029a", x"000030e866773ba7", 120539975, 62);
send(0, x"0000000000000265", x"00002d0fb54f8023", 40297172, 62);
send(1, x"0000000000000199", x"000037646a86cff1", -80509018, 62);
send(2, x"0000000000000295", x"000033affbdfdcdd", 161337941, 62);
send(3, x"0000000000000259", x"000030e870a73c1a", 120539903, 62);
send(0, x"000000000000016a", x"00002d0fb40ab1db", 40297172, 62);
send(1, x"0000000000000156", x"0000376469a9a7bc", -80509018, 62);
send(2, x"0000000000000269", x"000033aff0ddacb7", 161337941, 62);
send(3, x"0000000000000256", x"000030e87ad74886", 120539903, 62);
send(0, x"00000000000002a5", x"00002d0fb2c5ec8f", 40297101, 62);
send(1, x"000000000000029a", x"0000376468cc8b82", -80509018, 62);
send(2, x"000000000000016a", x"000033afe5db7f8f", 161337941, 62);
send(3, x"0000000000000155", x"000030e885075aef", 120539903, 62);
send(0, x"000000000000031f", x"00002d0fb181333d", 40297101, 62);
send(1, x"000000000000031f", x"0000376467ef813e", -80509018, 62);
send(2, x"000000000000031f", x"000033afdad95b63", 161337941, 62);
send(3, x"000000000000031f", x"000030e88f377953", 120539903, 62);
send(0, x"00000000000000ae", x"00002d0fb03c85e5", 40297101, 62);
send(1, x"00000000000000ae", x"00003764671282f5", -80509018, 62);
send(2, x"00000000000000ae", x"000033afcfd73d34", 161337941, 62);
send(3, x"00000000000000ae", x"000030e89967a0b2", 120539903, 62);
send(0, x"00000000000001a4", x"00002d0faef7e487", 40297101, 62);
send(1, x"00000000000001a4", x"00003764663590a5", -80509018, 62);
send(2, x"00000000000001a4", x"000033afc4d52204", 161337941, 62);
send(3, x"00000000000001a4", x"000030e8a397d10d", 120539903, 62);
send(0, x"000000000000026a", x"00002d0fadb34c25", 40297101, 62);
send(1, x"000000000000026a", x"000037646558b34b", -80509018, 62);
send(2, x"000000000000026a", x"000033afb9d30fcf", 161337941, 62);
send(3, x"000000000000026a", x"000030e8adc80d61", 120539903, 62);
send(0, x"0000000000000155", x"00002d0fac6ebfbc", 40297101, 62);
send(1, x"0000000000000155", x"00003764647be1eb", -80509018, 62);
send(2, x"0000000000000155", x"000033afaed10397", 161337941, 62);
send(3, x"00000000000002a9", x"000030e8b7f852b1", 120539903, 62);
send(0, x"0000000000000155", x"00002d0fab2a3f4e", 40297101, 62);
send(1, x"0000000000000155", x"00003764639f1c85", -80509018, 62);
send(2, x"0000000000000155", x"000033afa3cefa5d", 161337941, 62);
send(3, x"00000000000002aa", x"000030e8c228a0fc", 120539903, 62);
send(0, x"00000000000002a9", x"00002d0fa9e5c7db", 40297101, 62);
send(1, x"0000000000000156", x"0000376462c26916", -80509018, 62);
send(2, x"0000000000000156", x"000033af98ccfa20", 161337941, 62);
send(3, x"0000000000000156", x"000030e8cc58f844", 120539903, 62);
send(0, x"000000000000016a", x"00002d0fa8a15c61", 40297101, 62);
send(1, x"0000000000000255", x"0000376461e5c1a1", -80509090, 62);
send(2, x"0000000000000155", x"000033af8dcaffdf", 161337941, 62);
send(3, x"0000000000000269", x"000030e8d6895b85", 120539903, 62);
send(0, x"00000000000001aa", x"00002d0fa75cfce2", 40297101, 62);
send(1, x"0000000000000165", x"0000376461092c23", -80509090, 62);
send(2, x"00000000000002a6", x"000033af82c90e99", 161337941, 62);
send(3, x"0000000000000155", x"000030e8e0b9c7c1", 120539903, 62);
send(0, x"00000000000001aa", x"00002d0fa618a361", 40297101, 62);
send(1, x"0000000000000199", x"00003764602c9fa0", -80509090, 62);
send(2, x"0000000000000199", x"000033af77c71d54", 161337941, 62);
send(3, x"0000000000000295", x"000030e8eaea3cf9", 120539903, 62);
send(0, x"0000000000000166", x"00002d0fa4d458d7", 40297101, 62);
send(1, x"0000000000000165", x"000037645f502813", -80509090, 62);
send(2, x"0000000000000196", x"000033af6cc53509", 161337941, 62);
send(3, x"00000000000002a9", x"000030e8f51abe2b", 120539903, 62);
send(0, x"0000000000000266", x"00002d0fa3901a48", 40297101, 62);
send(1, x"0000000000000195", x"000037645e73bc81", -80509090, 62);
send(2, x"0000000000000199", x"000033af61c352bd", 161337941, 62);
send(3, x"0000000000000295", x"000030e8ff4b455a", 120539903, 62);
send(0, x"000000000000016a", x"00002d0fa24be4b4", 40297101, 62);
send(1, x"000000000000026a", x"000037645d975ce8", -80509090, 62);
send(2, x"0000000000000155", x"000033af56c1766d", 161337941, 62);
send(3, x"000000000000016a", x"000030e9097bd883", 120539903, 62);
send(0, x"0000000000000265", x"00002d0fa107bb19", 40297101, 62);
send(1, x"0000000000000256", x"000037645cbb0f46", -80509090, 62);
send(2, x"0000000000000169", x"000033af4bbfa01a", 161337941, 62);
send(3, x"0000000000000295", x"000030e913ac74a8", 120539903, 62);
send(0, x"0000000000000159", x"00002d0f9fc39a7b", 40297101, 62);
send(1, x"00000000000001a9", x"000037645bded09c", -80509090, 62);
send(2, x"0000000000000266", x"000033af40bdd2c2", 161337869, 62);
send(3, x"0000000000000165", x"000030e91ddd1cc6", 120539903, 62);
send(0, x"0000000000000295", x"00002d0f9e7f88d5", 40297101, 62);
send(1, x"0000000000000295", x"000037645b029dec", -80509090, 62);
send(2, x"00000000000002aa", x"000033af35bc056b", 161337869, 62);
send(3, x"000000000000016a", x"000030e9280dcae2", 120539903, 62);
send(0, x"00000000000002a6", x"00002d0f9d3b802b", 40297029, 62);
send(1, x"0000000000000169", x"000037645a267a36", -80509090, 62);
send(2, x"00000000000002a5", x"000033af2aba440d", 161337869, 62);
send(3, x"00000000000001a5", x"000030e9323e84f7", 120539903, 62);
send(0, x"000000000000019a", x"00002d0f9bf7807c", 40297029, 62);
send(1, x"000000000000026a", x"00003764594a6876", -80509090, 62);
send(2, x"00000000000001a6", x"000033af1fb885ae", 161337869, 62);
send(3, x"00000000000002a6", x"000030e93c6f4808", 120539831, 62);
send(0, x"0000000000000255", x"00002d0f9ab38fc5", 40297029, 62);
send(1, x"00000000000001a9", x"00003764586e62af", -80509090, 62);
send(2, x"0000000000000266", x"000033af14b6d04b", 161337869, 62);
send(3, x"000000000000025a", x"000030e946a01a11", 120539831, 62);
send(0, x"0000000000000169", x"00002d0f996fa50c", 40297029, 62);
send(1, x"00000000000002a6", x"00003764579268e4", -80509090, 62);
send(2, x"0000000000000166", x"000033af09b51de6", 161337869, 62);
send(3, x"000000000000016a", x"000030e950d0ef1a", 120539831, 62);
send(0, x"000000000000031f", x"00002d0f982bc64c", 40297029, 62);
send(1, x"000000000000031f", x"0000376456b6810f", -80509161, 62);
send(2, x"000000000000031f", x"000033aefeb3717e", 161337869, 62);
send(3, x"000000000000031f", x"000030e95b01d01c", 120539831, 62);
send(0, x"00000000000000ae", x"00002d0f96e7f685", 40297029, 62);
send(1, x"00000000000000ae", x"0000376455daa832", -80509161, 62);
send(2, x"00000000000000ae", x"000033aef3b1ce11", 161337869, 62);
send(3, x"00000000000000ae", x"000030e96532ba19", 120539831, 62);
send(0, x"00000000000001a4", x"00002d0f95a42fba", 40297029, 62);
send(1, x"00000000000001a4", x"0000376454fedb50", -80509161, 62);
send(2, x"00000000000001a4", x"000033aee8b02da3", 161337869, 62);
send(3, x"00000000000001a4", x"000030e96f63b011", 120539831, 62);
send(0, x"000000000000015a", x"00002d0f946071e9", 40297029, 62);
send(1, x"000000000000015a", x"0000376454232064", -80509161, 62);
send(2, x"000000000000015a", x"000033aeddae9631", 161337869, 62);
send(3, x"000000000000015a", x"000030e97994ac05", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f931cc312", 40297029, 62);
send(1, x"00000000000001aa", x"0000376453477173", -80509161, 62);
send(2, x"00000000000002aa", x"000033aed2ad04bb", 161337869, 62);
send(3, x"0000000000000155", x"000030e983c5b3f3", 120539831, 62);
send(0, x"0000000000000195", x"00002d0f91d91d36", 40297029, 62);
send(1, x"0000000000000169", x"00003764526bd17a", -80509161, 62);
send(2, x"00000000000001a6", x"000033aec7ab7346", 161337869, 62);
send(3, x"00000000000002a6", x"000030e98df6c4de", 120539831, 62);
send(0, x"0000000000000199", x"00002d0f90958056", 40297029, 62);
send(1, x"00000000000001a6", x"0000376451904079", -80509161, 62);
send(2, x"0000000000000299", x"000033aebca9edca", 161337869, 62);
send(3, x"00000000000001a6", x"000030e99827e1c2", 120539831, 62);
send(0, x"0000000000000255", x"00002d0f8f51ef6f", 40297029, 62);
send(1, x"0000000000000269", x"0000376450b4be71", -80509161, 62);
send(2, x"000000000000026a", x"000033aeb1a86e4b", 161337869, 62);
send(3, x"000000000000029a", x"000030e9a25907a1", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f8e0e6a83", 40297029, 62);
send(1, x"0000000000000156", x"000037644fd94b62", -80509161, 62);
send(2, x"00000000000002aa", x"000033aea6a6f4ca", 161337869, 62);
send(3, x"00000000000002a9", x"000030e9ac8a367c", 120539831, 62);
send(0, x"00000000000001aa", x"00002d0f8ccaee91", 40297029, 62);
send(1, x"0000000000000255", x"000037644efde44c", -80509161, 62);
send(2, x"00000000000001aa", x"000033ae9ba57e47", 161337869, 62);
send(3, x"00000000000001aa", x"000030e9b6bb7151", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f8b877e9a", 40297029, 62);
send(1, x"0000000000000155", x"000037644e228f2e", -80509161, 62);
send(2, x"00000000000002aa", x"000033ae90a413be", 161337869, 62);
send(3, x"00000000000002aa", x"000030e9c0ecb223", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f8a441a9e", 40297029, 62);
send(1, x"0000000000000155", x"000037644d474908", -80509161, 62);
send(2, x"00000000000002aa", x"000033ae85a2ac33", 161337869, 62);
send(3, x"00000000000002aa", x"000030e9cb1dfeef", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f8900c29a", 40297029, 62);
send(1, x"0000000000000155", x"000037644c6c0bdd", -80509161, 62);
send(2, x"00000000000002aa", x"000033ae7aa147a8", 161337869, 62);
send(3, x"00000000000002aa", x"000030e9d54f54b6", 120539831, 62);
send(0, x"00000000000001a6", x"00002d0f87bd7393", 40296957, 62);
send(1, x"0000000000000259", x"000037644b90e3a8", -80509233, 62);
send(2, x"00000000000001a6", x"000033ae6f9fec17", 161337869, 62);
send(3, x"00000000000001a6", x"000030e9df80b37a", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f867a3086", 40296957, 62);
send(1, x"0000000000000155", x"000037644ab5c76d", -80509233, 62);
send(2, x"00000000000002aa", x"000033ae649e9684", 161337869, 62);
send(3, x"00000000000002aa", x"000030e9e9b21b38", 120539831, 62);
send(0, x"00000000000002aa", x"00002d0f8536f972", 40296957, 62);
send(1, x"0000000000000155", x"0000376449dab72c", -80509233, 62);
send(2, x"00000000000002aa", x"000033ae599d46ed", 161337869, 62);
send(3, x"00000000000002aa", x"000030e9f3e38ef1", 120539831, 62);
send(0, x"00000000000002a6", x"00002d0f83f3cb5a", 40296957, 62);
send(1, x"0000000000000159", x"0000376448ffb8e2", -80509233, 62);
send(2, x"00000000000002a6", x"000033ae4e9bfd54", 161337869, 62);
send(3, x"00000000000002a6", x"000030e9fe150ba5", 120539760, 62);
send(0, x"00000000000001aa", x"00002d0f82b0a93c", 40296957, 62);
send(1, x"000000000000016a", x"000037644824c991", -80509233, 62);
send(2, x"000000000000015a", x"000033ae439ab9b7", 161337869, 62);
send(3, x"000000000000026a", x"000030ea08469154", 120539760, 62);
send(0, x"00000000000001a5", x"00002d0f816d9318", 40296957, 62);
send(1, x"0000000000000165", x"000037644749e937", -80509233, 62);
send(2, x"0000000000000165", x"000033ae38997f16", 161337869, 62);
send(3, x"000000000000026a", x"000030ea127825fc", 120539760, 62);
send(0, x"000000000000016a", x"00002d0f802a82f1", 40296957, 62);
send(1, x"00000000000002aa", x"00003764466f14d8", -80509233, 62);
send(2, x"0000000000000295", x"000033ae2d984475", 161337869, 62);
send(3, x"0000000000000156", x"000030ea1ca9c0a1", 120539760, 62);
send(0, x"000000000000031f", x"00002d0f7ee781c2", 40296957, 62);
send(1, x"000000000000031f", x"0000376445944f72", -80509233, 62);
send(2, x"000000000000031f", x"000033ae229715ce", 161337869, 62);
send(3, x"000000000000031f", x"000030ea26db6442", 120539760, 62);
send(0, x"00000000000000ae", x"00002d0f7da48c8e", 40296957, 62);
send(1, x"00000000000000ae", x"0000376444b99c03", -80509233, 62);
send(2, x"00000000000000ae", x"000033ae1795ea26", 161337869, 62);
send(3, x"00000000000000ae", x"000030ea310d10de", 120539760, 62);
send(0, x"00000000000001a4", x"00002d0f7c61a055", 40296957, 62);
send(1, x"00000000000001a4", x"0000376443def18e", -80509233, 62);
send(2, x"00000000000001a4", x"000033ae0c94c47a", 161337869, 62);
send(3, x"00000000000001a4", x"000030ea3b3ec675", 120539760, 62);
send(0, x"000000000000025a", x"00002d0f7b1ec016", 40296957, 62);
send(1, x"000000000000025a", x"0000376443045911", -80509233, 62);
send(2, x"000000000000025a", x"000033ae0193a7ca", 161337869, 62);
send(3, x"000000000000025a", x"000030ea45708806", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f79dbebd1", 40296957, 62);
send(1, x"00000000000002aa", x"000037644229cf8d", -80509233, 62);
send(2, x"00000000000002aa", x"000033adf6928e19", 161337869, 62);
send(3, x"00000000000002aa", x"000030ea4fa25294", 120539760, 62);
send(0, x"000000000000029a", x"00002d0f78992088", 40296957, 62);
send(1, x"000000000000029a", x"00003764414f5203", -80509233, 62);
send(2, x"000000000000029a", x"000033adeb917a64", 161337797, 62);
send(3, x"000000000000029a", x"000030ea59d4291b", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f77566138", 40296957, 62);
send(1, x"00000000000002aa", x"000037644074e66f", -80509305, 62);
send(2, x"00000000000002aa", x"000033ade0906fab", 161337797, 62);
send(3, x"00000000000002aa", x"000030ea6406059f", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f7613ade3", 40296957, 62);
send(1, x"00000000000002aa", x"000037643f9a89d4", -80509305, 62);
send(2, x"00000000000002aa", x"000033add58f6aef", 161337797, 62);
send(3, x"00000000000002aa", x"000030ea6e37ee1d", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f74d10389", 40296957, 62);
send(1, x"00000000000002aa", x"000037643ec03933", -80509305, 62);
send(2, x"00000000000002aa", x"000033adca8e6932", 161337797, 62);
send(3, x"00000000000002aa", x"000030ea7869e294", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f738e622a", 40296957, 62);
send(1, x"00000000000002aa", x"000037643de5f78b", -80509305, 62);
send(2, x"00000000000002aa", x"000033adbf8d6d71", 161337797, 62);
send(3, x"00000000000002aa", x"000030ea829bdd0a", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f724bcfc4", 40296886, 62);
send(1, x"00000000000002aa", x"000037643d0bc4db", -80509305, 62);
send(2, x"00000000000002aa", x"000033adb48c7aac", 161337797, 62);
send(3, x"00000000000002aa", x"000030ea8ccde379", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f7109465a", 40296886, 62);
send(1, x"00000000000002aa", x"000037643c31a123", -80509305, 62);
send(2, x"00000000000002aa", x"000033ada98b8de4", 161337797, 62);
send(3, x"00000000000002aa", x"000030ea96fff2e3", 120539760, 62);
send(0, x"00000000000002aa", x"00002d0f6fc6c8e9", 40296886, 62);
send(1, x"00000000000002aa", x"000037643b578966", -80509305, 62);
send(2, x"00000000000002aa", x"000033ad9e8aa41b", 161337797, 62);
send(3, x"00000000000002aa", x"000030eaa1320b49", 120539760, 62);
send(0, x"0000000000000166", x"00002d0f6e845773", 40296886, 62);
send(1, x"0000000000000166", x"000037643a7d839f", -80509305, 62);
send(2, x"0000000000000166", x"000033ad9389c34d", 161337797, 62);
send(3, x"0000000000000166", x"000030eaab642cab", 120539760, 62);
send(0, x"0000000000000155", x"00002d0f6d41eef8", 40296886, 62);
send(1, x"0000000000000155", x"0000376439a38cd1", -80509305, 62);
send(2, x"0000000000000155", x"000033ad8888e87c", 161337797, 62);
send(3, x"0000000000000155", x"000030eab5965a06", 120539760, 62);
send(0, x"0000000000000155", x"00002d0f6bff9277", 40296886, 62);
send(1, x"0000000000000155", x"0000376438c9a1fd", -80509305, 62);
send(2, x"0000000000000155", x"000033ad7d8813a8", 161337797, 62);
send(3, x"0000000000000155", x"000030eabfc88d5f", 120539688, 62);
send(0, x"0000000000000155", x"00002d0f6abd41f0", 40296886, 62);
send(1, x"0000000000000155", x"0000376437efc622", -80509305, 62);
send(2, x"0000000000000155", x"000033ad728744d1", 161337797, 62);
send(3, x"0000000000000155", x"000030eac9faccb1", 120539688, 62);
send(0, x"0000000000000155", x"00002d0f697afa64", 40296886, 62);
send(1, x"0000000000000155", x"000037643715fc3d", -80509305, 62);
send(2, x"0000000000000155", x"000033ad67867bf7", 161337797, 62);
send(3, x"0000000000000155", x"000030ead42d17fe", 120539688, 62);
send(0, x"0000000000000155", x"00002d0f6838bed3", 40296886, 62);
send(1, x"0000000000000155", x"00003764363c3e53", -80509305, 62);
send(2, x"0000000000000155", x"000033ad5c85b919", 161337797, 62);
send(3, x"0000000000000155", x"000030eade5f6c46", 120539688, 62);
send(0, x"0000000000000159", x"00002d0f66f68c3d", 40296886, 62);
send(1, x"0000000000000159", x"0000376435628c62", -80509376, 62);
send(2, x"0000000000000159", x"000033ad5184fc39", 161337797, 62);
send(3, x"0000000000000159", x"000030eae891c989", 120539688, 62);
send(0, x"000000000000031f", x"00002d0f65b465a1", 40296886, 62);
send(1, x"000000000000031f", x"000037643488ec69", -80509376, 62);
send(2, x"000000000000031f", x"000033ad46844557", 161337797, 62);
send(3, x"000000000000031f", x"000030eaf2c42fc8", 120539688, 62);
send(0, x"00000000000000ae", x"00002d0f64724aff", 40296886, 62);
send(1, x"00000000000000ae", x"0000376433af5b67", -80509376, 62);
send(2, x"00000000000000ae", x"000033ad3b839471", 161337797, 62);
send(3, x"00000000000000ae", x"000030eafcf6a201", 120539688, 62);
send(0, x"00000000000001a4", x"00002d0f63303c57", 40296886, 62);
send(1, x"00000000000001a4", x"0000376432d5d661", -80509376, 62);
send(2, x"00000000000001a4", x"000033ad3082e987", 161337797, 62);
send(3, x"00000000000001a4", x"000030eb07291a37", 120539688, 62);
send(0, x"000000000000029a", x"00002d0f61ee36aa", 40296886, 62);
send(1, x"000000000000029a", x"0000376431fc6052", -80509376, 62);
send(2, x"000000000000029a", x"000033ad2582449c", 161337797, 62);
send(3, x"000000000000029a", x"000030eb115b9e67", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f60ac3cf8", 40296886, 62);
send(1, x"00000000000002aa", x"000037643122fc3b", -80509376, 62);
send(2, x"00000000000002aa", x"000033ad1a81a8ab", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb1b8e2b93", 120539688, 62);
send(0, x"000000000000029a", x"00002d0f5f6a4f3f", 40296886, 62);
send(1, x"000000000000029a", x"000037643049a11f", -80509376, 62);
send(2, x"000000000000029a", x"000033ad0f810fb9", 161337797, 62);
send(3, x"000000000000029a", x"000030eb25c0c4b8", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f5e286a82", 40296886, 62);
send(1, x"00000000000002aa", x"000037642f705af8", -80509376, 62);
send(2, x"00000000000002aa", x"000033ad04807cc4", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb2ff363db", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f5ce691bf", 40296814, 62);
send(1, x"00000000000002aa", x"000037642e9720cc", -80509376, 62);
send(2, x"00000000000002aa", x"000033acf97ff2ca", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb3a260ef7", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f5ba4c4f6", 40296814, 62);
send(1, x"00000000000002aa", x"000037642dbdf598", -80509376, 62);
send(2, x"00000000000002aa", x"000033acee7f6ece", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb4458c60e", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f5a62fe2a", 40296814, 62);
send(1, x"00000000000002aa", x"000037642ce4d65e", -80509376, 62);
send(2, x"00000000000002aa", x"000033ace37eead2", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb4e8b8321", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f59214657", 40296814, 62);
send(1, x"00000000000002aa", x"000037642c0bc91a", -80509376, 62);
send(2, x"00000000000002aa", x"000033acd87e72cf", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb58be4c2f", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f57df9a7d", 40296814, 62);
send(1, x"00000000000002aa", x"000037642b32c7d2", -80509448, 62);
send(2, x"00000000000002aa", x"000033accd7e00c9", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb62f11e38", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f569df79f", 40296814, 62);
send(1, x"00000000000002aa", x"000037642a59d581", -80509448, 62);
send(2, x"00000000000002aa", x"000033acc27d91c3", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb6d23f93c", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f555c60bb", 40296814, 62);
send(1, x"00000000000002aa", x"000037642980f229", -80509448, 62);
send(2, x"00000000000002aa", x"000033acb77d2bb7", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb7756e03b", 120539688, 62);
send(0, x"00000000000002aa", x"00002d0f541ad5d1", 40296814, 62);
send(1, x"00000000000002aa", x"0000376428a81dca", -80509448, 62);
send(2, x"00000000000002aa", x"000033acac7ccba9", 161337797, 62);
send(3, x"00000000000002aa", x"000030eb8189cd36", 120539617, 62);
send(0, x"00000000000002aa", x"00002d0f52d953e3", 40296814, 62);
send(1, x"00000000000002aa", x"0000376427cf5862", -80509448, 62);
send(2, x"00000000000002aa", x"000033aca17c6e99", 161337726, 62);
send(3, x"00000000000002aa", x"000030eb8bbcc62c", 120539617, 62);
send(0, x"00000000000002aa", x"00002d0f5197ddee", 40296814, 62);
send(1, x"00000000000002aa", x"0000376426f6a1f4", -80509448, 62);
send(2, x"00000000000002aa", x"000033ac967c1a84", 161337726, 62);
send(3, x"00000000000002aa", x"000030eb95efc81c", 120539617, 62);
send(0, x"00000000000002aa", x"00002d0f505673f4", 40296814, 62);
send(1, x"00000000000002aa", x"00003764261dfa7e", -80509448, 62);
send(2, x"00000000000002aa", x"000033ac8b7bcc6d", 161337726, 62);
send(3, x"00000000000002aa", x"000030eba022d607", 120539617, 62);
send(0, x"00000000000001aa", x"00002d0f4f1512f5", 40296814, 62);
send(1, x"00000000000001aa", x"0000376425455f02", -80509448, 62);
send(2, x"00000000000001aa", x"000033ac807b8452", 161337726, 62);
send(3, x"00000000000001aa", x"000030ebaa55ecee", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f4dd3baf1", 40296814, 62);
send(1, x"0000000000000155", x"00003764246cd27f", -80509448, 62);
send(2, x"0000000000000155", x"000033ac757b4235", 161337726, 62);
send(3, x"0000000000000155", x"000030ebb4890cd0", 120539617, 62);
send(0, x"000000000000031f", x"00002d0f4c9271e6", 40296814, 62);
send(1, x"000000000000031f", x"00003764239457f2", -80509448, 62);
send(2, x"000000000000031f", x"000033ac6a7b0614", 161337726, 62);
send(3, x"000000000000031f", x"000030ebbebc35ae", 120539617, 62);
send(0, x"00000000000000ae", x"00002d0f4b5131d7", 40296814, 62);
send(1, x"00000000000000ae", x"0000376422bbe960", -80509448, 62);
send(2, x"00000000000000ae", x"000033ac5f7acff0", 161337726, 62);
send(3, x"00000000000000ae", x"000030ebc8ef6a85", 120539617, 62);
send(0, x"00000000000001a4", x"00002d0f4a0ffdc1", 40296814, 62);
send(1, x"00000000000001a4", x"0000376421e386c7", -80509448, 62);
send(2, x"00000000000001a4", x"000033ac547a9fca", 161337726, 62);
send(3, x"00000000000001a4", x"000030ebd322a55a", 120539617, 62);
send(0, x"000000000000019a", x"00002d0f48ced5a6", 40296814, 62);
send(1, x"000000000000019a", x"00003764210b3626", -80509448, 62);
send(2, x"000000000000019a", x"000033ac497a75a1", 161337726, 62);
send(3, x"000000000000019a", x"000030ebdd55ec28", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f478db686", 40296743, 62);
send(1, x"0000000000000155", x"000037642032f47c", -80509519, 62);
send(2, x"0000000000000155", x"000033ac3e7a5174", 161337726, 62);
send(3, x"0000000000000155", x"000030ebe7893bf2", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f464ca360", 40296743, 62);
send(1, x"0000000000000155", x"000037641f5abece", -80509519, 62);
send(2, x"0000000000000155", x"000033ac337a3345", 161337726, 62);
send(3, x"0000000000000155", x"000030ebf1bc97b6", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f450b9c34", 40296743, 62);
send(1, x"0000000000000155", x"000037641e829b15", -80509519, 62);
send(2, x"0000000000000155", x"000033ac287a1b12", 161337726, 62);
send(3, x"0000000000000155", x"000030ebfbeffc76", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f43ca9e03", 40296743, 62);
send(1, x"0000000000000155", x"000037641daa8656", -80509519, 62);
send(2, x"0000000000000155", x"000033ac1d7a0bdb", 161337726, 62);
send(3, x"0000000000000155", x"000030ec06236732", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f4289abcc", 40296743, 62);
send(1, x"0000000000000155", x"000037641cd27d91", -80509519, 62);
send(2, x"0000000000000155", x"000033ac127a02a1", 161337726, 62);
send(3, x"0000000000000155", x"000030ec1056e3e6", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f4148c292", 40296743, 62);
send(1, x"0000000000000155", x"000037641bfa83c3", -80509519, 62);
send(2, x"0000000000000155", x"000033ac0779f967", 161337726, 62);
send(3, x"0000000000000155", x"000030ec1a8a6398", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f4007e551", 40296743, 62);
send(1, x"0000000000000155", x"000037641b2298ef", -80509519, 62);
send(2, x"0000000000000155", x"000033abfc79fc27", 161337726, 62);
send(3, x"0000000000000155", x"000030ec24bdef44", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f3ec7140a", 40296743, 62);
send(1, x"0000000000000155", x"000037641a4abd13", -80509519, 62);
send(2, x"0000000000000155", x"000033abf17a04e4", 161337726, 62);
send(3, x"0000000000000155", x"000030ec2ef183eb", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f3d864bbe", 40296743, 62);
send(1, x"0000000000000155", x"000037641972ed31", -80509519, 62);
send(2, x"0000000000000155", x"000033abe67a10a0", 161337726, 62);
send(3, x"0000000000000155", x"000030ec3925218e", 120539617, 62);
send(0, x"0000000000000155", x"00002d0f3c45926b", 40296743, 62);
send(1, x"0000000000000155", x"00003764189b2f46", -80509519, 62);
send(2, x"0000000000000155", x"000033abdb7a2556", 161337726, 62);
send(3, x"0000000000000155", x"000030ec4358c82d", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f3b04e214", 40296743, 62);
send(1, x"0000000000000155", x"0000376417c38054", -80509519, 62);
send(2, x"0000000000000155", x"000033abd07a3d0c", 161337726, 62);
send(3, x"0000000000000155", x"000030ec4d8c7ac5", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f39c43ab8", 40296743, 62);
send(1, x"0000000000000155", x"0000376416ebdd5b", -80509519, 62);
send(2, x"0000000000000155", x"000033abc57a5abf", 161337726, 62);
send(3, x"0000000000000155", x"000030ec57c03659", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f3883a254", 40296743, 62);
send(1, x"0000000000000155", x"000037641614495b", -80509519, 62);
send(2, x"0000000000000155", x"000033abba7a816c", 161337726, 62);
send(3, x"0000000000000155", x"000030ec61f3fae9", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f374312ec", 40296743, 62);
send(1, x"0000000000000155", x"00003764153cc752", -80509591, 62);
send(2, x"0000000000000155", x"000033abaf7aae18", 161337726, 62);
send(3, x"0000000000000155", x"000030ec6c27c873", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f36028c80", 40296743, 62);
send(1, x"0000000000000155", x"0000376414655143", -80509591, 62);
send(2, x"0000000000000155", x"000033aba47ae3be", 161337726, 62);
send(3, x"0000000000000155", x"000030ec765ba4f7", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f34c2120d", 40296743, 62);
send(1, x"0000000000000155", x"00003764138de72e", -80509591, 62);
send(2, x"0000000000000155", x"000033ab997b1964", 161337726, 62);
send(3, x"0000000000000155", x"000030ec808f8777", 120539545, 62);
send(0, x"000000000000031f", x"00002d0f3381a395", 40296743, 62);
send(1, x"000000000000031f", x"0000376412b68f10", -80509591, 62);
send(2, x"000000000000031f", x"000033ab8e7b5807", 161337726, 62);
send(3, x"000000000000031f", x"000030ec8ac372f4", 120539545, 62);
send(0, x"00000000000000ae", x"00002d0f32413e18", 40296671, 62);
send(1, x"00000000000000ae", x"0000376411df45ea", -80509591, 62);
send(2, x"00000000000000ae", x"000033ab837b9ca5", 161337726, 62);
send(3, x"00000000000000ae", x"000030ec94f76a6a", 120539545, 62);
send(0, x"00000000000001a4", x"00002d0f3100e793", 40296671, 62);
send(1, x"00000000000001a4", x"00003764110808bf", -80509591, 62);
send(2, x"00000000000001a4", x"000033ab787be443", 161337726, 62);
send(3, x"00000000000001a4", x"000030ec9f2b67dd", 120539545, 62);
send(0, x"0000000000000156", x"00002d0f2fc0970c", 40296671, 62);
send(1, x"0000000000000156", x"000037641030da8c", -80509591, 62);
send(2, x"0000000000000156", x"000033ab6d7c37db", 161337726, 62);
send(3, x"0000000000000156", x"000030eca95f7149", 120539545, 62);
send(0, x"0000000000000295", x"00002d0f2e80557d", 40296671, 62);
send(1, x"0000000000000295", x"000037640f59be50", -80509591, 62);
send(2, x"0000000000000295", x"000033ab627c8e71", 161337726, 62);
send(3, x"0000000000000295", x"000030ecb39386b1", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f2d401ce9", 40296671, 62);
send(1, x"0000000000000155", x"000037640e82ab10", -80509591, 62);
send(2, x"0000000000000155", x"000033ab577ceb04", 161337726, 62);
send(3, x"0000000000000155", x"000030ecbdc7a215", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f2bfff050", 40296671, 62);
send(1, x"0000000000000155", x"000037640dabacc4", -80509591, 62);
send(2, x"0000000000000155", x"000033ab4c7d4d94", 161337654, 62);
send(3, x"0000000000000155", x"000030ecc7fbc972", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f2abfcfb0", 40296671, 62);
send(1, x"0000000000000155", x"000037640cd4ba74", -80509591, 62);
send(2, x"0000000000000155", x"000033ab417db91f", 161337654, 62);
send(3, x"0000000000000155", x"000030ecd22ff9cc", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f297fb80c", 40296671, 62);
send(1, x"0000000000000155", x"000037640bfdd71b", -80509591, 62);
send(2, x"0000000000000155", x"000033ab367e27a9", 161337654, 62);
send(3, x"0000000000000155", x"000030ecdc643620", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f283fa963", 40296671, 62);
send(1, x"0000000000000155", x"000037640b26ffbd", -80509591, 62);
send(2, x"0000000000000155", x"000033ab2b7e9c30", 161337654, 62);
send(3, x"0000000000000155", x"000030ece6987870", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f26ffa9b4", 40296671, 62);
send(1, x"0000000000000155", x"000037640a503a55", -80509663, 62);
send(2, x"0000000000000155", x"000033ab207f19b3", 161337654, 62);
send(3, x"0000000000000155", x"000030ecf0ccc6bb", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f25bfb2ff", 40296671, 62);
send(1, x"0000000000000155", x"00003764097980e8", -80509663, 62);
send(2, x"0000000000000155", x"000033ab157f9a34", 161337654, 62);
send(3, x"0000000000000155", x"000030ecfb011e01", 120539545, 62);
send(0, x"0000000000000155", x"00002d0f247fc845", 40296671, 62);
send(1, x"0000000000000155", x"0000376408a2d673", -80509663, 62);
send(2, x"0000000000000155", x"000033ab0a8020b2", 161337654, 62);
send(3, x"0000000000000155", x"000030ed05357e42", 120539474, 62);
send(0, x"0000000000000155", x"00002d0f233fe984", 40296671, 62);
send(1, x"0000000000000155", x"0000376407cc3af6", -80509663, 62);
send(2, x"0000000000000155", x"000033aaff80b02b", 161337654, 62);
send(3, x"0000000000000155", x"000030ed0f69e77f", 120539474, 62);
send(0, x"0000000000000155", x"00002d0f220013bf", 40296671, 62);
send(1, x"0000000000000155", x"0000376406f5ae72", -80509663, 62);
send(2, x"0000000000000155", x"000033aaf48145a1", 161337654, 62);
send(3, x"0000000000000155", x"000030ed199e5cb6", 120539474, 62);
send(0, x"0000000000000155", x"00002d0f20c049f4", 40296671, 62);
send(1, x"0000000000000155", x"00003764061f30e6", -80509663, 62);
send(2, x"0000000000000155", x"000033aae981de17", 161337654, 62);
send(3, x"0000000000000155", x"000030ed23d2dae9", 120539474, 62);
send(0, x"0000000000000155", x"00002d0f1f808c23", 40296671, 62);
send(1, x"0000000000000155", x"000037640548c254", -80509663, 62);
send(2, x"0000000000000155", x"000033aade827f87", 161337654, 62);
send(3, x"0000000000000155", x"000030ed2e076216", 120539474, 62);
send(0, x"0000000000000155", x"00002d0f1e40d74e", 40296671, 62);
send(1, x"0000000000000155", x"00003764047262b9", -80509663, 62);
send(2, x"0000000000000155", x"000033aad38326f4", 161337654, 62);
send(3, x"0000000000000155", x"000030ed383bf53f", 120539474, 62);
send(0, x"0000000000000195", x"00002d0f1d012e72", 40296600, 62);
send(1, x"0000000000000195", x"00003764039c0f19", -80509663, 62);
send(2, x"0000000000000195", x"000033aac883d45f", 161337654, 62);
send(3, x"0000000000000195", x"000030ed42709162", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f1bc18b93", 40296600, 62);
send(1, x"00000000000002aa", x"0000376402c5ca71", -80509663, 62);
send(2, x"00000000000002aa", x"000033aabd8484c8", 161337654, 62);
send(3, x"00000000000002aa", x"000030ed4ca53681", 120539474, 62);
send(0, x"000000000000031f", x"00002d0f1a81faac", 40296600, 62);
send(1, x"000000000000031f", x"0000376401ef97bf", -80509663, 62);
send(2, x"000000000000031f", x"000033aab2853e2d", 161337654, 62);
send(3, x"000000000000031f", x"000030ed56d9e79a", 120539474, 62);
send(0, x"00000000000000ae", x"00002d0f194272c0", 40296600, 62);
send(1, x"00000000000000ae", x"0000376401197108", -80509663, 62);
send(2, x"00000000000000ae", x"000033aaa785fd8e", 161337654, 62);
send(3, x"00000000000000ae", x"000030ed610e9eb0", 120539474, 62);
send(0, x"00000000000001a4", x"00002d0f1802f3d0", 40296600, 62);
send(1, x"00000000000001a4", x"000037640043564c", -80509663, 62);
send(2, x"00000000000001a4", x"000033aa9c86bfee", 161337654, 62);
send(3, x"00000000000001a4", x"000030ed6b4361c0", 120539474, 62);
send(0, x"0000000000000256", x"00002d0f16c383d8", 40296600, 62);
send(1, x"0000000000000256", x"00003763ff6d4d86", -80509734, 62);
send(2, x"0000000000000256", x"000033aa91878e48", 161337654, 62);
send(3, x"0000000000000256", x"000030ed75782dcc", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f15841cdb", 40296600, 62);
send(1, x"00000000000002aa", x"00003763fe9753b8", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa86885fa1", 161337654, 62);
send(3, x"00000000000002aa", x"000030ed7fad02d3", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f1444beda", 40296600, 62);
send(1, x"00000000000002aa", x"00003763fdc165e5", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa7b8936f6", 161337654, 62);
send(3, x"00000000000002aa", x"000030ed89e1e0d5", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f13056cd3", 40296600, 62);
send(1, x"00000000000002aa", x"00003763fceb8a08", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa708a1449", 161337654, 62);
send(3, x"00000000000002aa", x"000030ed9416cad1", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f11c626c6", 40296600, 62);
send(1, x"00000000000002aa", x"00003763fc15bd24", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa658af798", 161337654, 62);
send(3, x"00000000000002aa", x"000030ed9e4bbdc9", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f1086ecb3", 40296600, 62);
send(1, x"00000000000002aa", x"00003763fb3ffc3a", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa5a8be3e3", 161337654, 62);
send(3, x"00000000000002aa", x"000030eda880bcbc", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f0f47b89d", 40296600, 62);
send(1, x"00000000000002aa", x"00003763fa6a4a48", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa4f8cd32d", 161337654, 62);
send(3, x"00000000000002aa", x"000030edb2b5c1ab", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f0e08937f", 40296600, 62);
send(1, x"00000000000002aa", x"00003763f994a750", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa448dc873", 161337654, 62);
send(3, x"00000000000002aa", x"000030edbcead294", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f0cc97a5c", 40296600, 62);
send(1, x"00000000000002aa", x"00003763f8bf134f", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa398ec6b5", 161337654, 62);
send(3, x"00000000000002aa", x"000030edc71fec78", 120539474, 62);
send(0, x"00000000000002aa", x"00002d0f0b8a6a34", 40296600, 62);
send(1, x"00000000000002aa", x"00003763f7e98b49", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa2e8fc7f5", 161337654, 62);
send(3, x"00000000000002aa", x"000030edd1550f58", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0f0a4b6606", 40296600, 62);
send(1, x"00000000000002aa", x"00003763f7141539", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa2390d232", 161337654, 62);
send(3, x"00000000000002aa", x"000030eddb8a3e32", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0f090c6ad3", 40296600, 62);
send(1, x"00000000000002aa", x"00003763f63eae22", -80509734, 62);
send(2, x"00000000000002aa", x"000033aa1891df6c", 161337654, 62);
send(3, x"00000000000002aa", x"000030ede5bf7309", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0f07cd7e99", 40296528, 62);
send(1, x"00000000000002aa", x"00003763f5695305", -80509806, 62);
send(2, x"00000000000002aa", x"000033aa0d92f2a3", 161337654, 62);
send(3, x"00000000000002aa", x"000030edeff4b3da", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0f068e9b5b", 40296528, 62);
send(1, x"00000000000002aa", x"00003763f49406e0", -80509806, 62);
send(2, x"00000000000002aa", x"000033aa02940ed7", 161337583, 62);
send(3, x"00000000000002aa", x"000030edfa29fda6", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0f054fc118", 40296528, 62);
send(1, x"00000000000002aa", x"00003763f3beccb3", -80509806, 62);
send(2, x"00000000000002aa", x"000033a9f7953106", 161337583, 62);
send(3, x"00000000000002aa", x"000030ee045f536d", 120539402, 62);
send(0, x"000000000000029a", x"00002d0f0410f2cf", 40296528, 62);
send(1, x"000000000000029a", x"00003763f2e99e80", -80509806, 62);
send(2, x"000000000000029a", x"000033a9ec965934", 161337583, 62);
send(3, x"000000000000029a", x"000030ee0e94b22f", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0f02d22d82", 40296528, 62);
send(1, x"00000000000002aa", x"00003763f2147c46", -80509806, 62);
send(2, x"00000000000002aa", x"000033a9e197875d", 161337583, 62);
send(3, x"00000000000002aa", x"000030ee18ca19ec", 120539402, 62);
send(0, x"000000000000031f", x"00002d0f0193772d", 40296528, 62);
send(1, x"000000000000031f", x"00003763f13f6c03", -80509806, 62);
send(2, x"000000000000031f", x"000033a9d698bb85", 161337583, 62);
send(3, x"000000000000031f", x"000030ee22ff8da4", 120539402, 62);
send(0, x"00000000000000ae", x"00002d0f0054c9d3", 40296528, 62);
send(1, x"00000000000000ae", x"00003763f06a6ab9", -80509806, 62);
send(2, x"00000000000000ae", x"000033a9cb99f5a9", 161337583, 62);
send(3, x"00000000000000ae", x"000030ee2d350759", 120539402, 62);
send(0, x"00000000000001a4", x"00002d0eff162874", 40296528, 62);
send(1, x"00000000000001a4", x"00003763ef957569", -80509806, 62);
send(2, x"00000000000001a4", x"000033a9c09b32cb", 161337583, 62);
send(3, x"00000000000001a4", x"000030ee376a8d07", 120539402, 62);
send(0, x"0000000000000296", x"00002d0efdd7930e", 40296528, 62);
send(1, x"0000000000000296", x"00003763eec09211", -80509806, 62);
send(2, x"0000000000000296", x"000033a9b59c7be8", 161337583, 62);
send(3, x"0000000000000296", x"000030ee41a01bb1", 120539402, 62);
send(0, x"00000000000002aa", x"00002d0efc9906a4", 40296528, 62);
send(1, x"00000000000002aa", x"00003763edebbab2", -80509806, 62);
send(2, x"00000000000002aa", x"000033a9aa9dc803", 161337583, 62);
send(3, x"00000000000002aa", x"000030ee4bd5b356", 120539402, 62);
send(0, x"0000000000000165", x"00002d0efb5a8634", 40296528, 62);
send(1, x"0000000000000165", x"00003763ed16f24b", -80509806, 62);
send(2, x"0000000000000165", x"000033a99f9f171c", 161337583, 62);
send(3, x"0000000000000165", x"000030ee560b53f8", 120539402, 62);
send(0, x"0000000000000155", x"00002d0efa1c0ec0", 40296528, 62);
send(1, x"0000000000000155", x"00003763ec4238dd", -80509806, 62);
send(2, x"0000000000000155", x"000033a994a07230", 161337583, 62);
send(3, x"0000000000000155", x"000030ee60410093", 120539402, 62);
send(0, x"0000000000000155", x"00002d0ef8dda644", 40296528, 62);
send(1, x"0000000000000155", x"00003763eb6d8e68", -80509806, 62);
send(2, x"0000000000000155", x"000033a989a1d041", 161337583, 62);
send(3, x"0000000000000155", x"000030ee6a76b629", 120539402, 62);
send(0, x"0000000000000155", x"00002d0ef79f43c5", 40296528, 62);
send(1, x"0000000000000155", x"00003763ea98f2eb", -80509877, 62);
send(2, x"0000000000000155", x"000033a97ea3374f", 161337583, 62);
send(3, x"0000000000000155", x"000030ee74ac77ba", 120539402, 62);
send(0, x"0000000000000155", x"00002d0ef660ed40", 40296528, 62);
send(1, x"0000000000000155", x"00003763e9c46367", -80509877, 62);
send(2, x"0000000000000155", x"000033a973a4a15b", 161337583, 62);
send(3, x"0000000000000155", x"000030ee7ee23f47", 120539402, 62);
send(0, x"0000000000000155", x"00002d0ef522a2b5", 40296528, 62);
send(1, x"0000000000000155", x"00003763e8efe5db", -80509877, 62);
send(2, x"0000000000000155", x"000033a968a61164", 161337583, 62);
send(3, x"0000000000000155", x"000030ee891812cf", 120539402, 62);
send(0, x"0000000000000155", x"00002d0ef3e46424", 40296528, 62);
send(1, x"0000000000000155", x"00003763e81b7748", -80509877, 62);
send(2, x"0000000000000155", x"000033a95da78a69", 161337583, 62);
send(3, x"0000000000000155", x"000030ee934def52", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ef2a6318d", 40296456, 62);
send(1, x"0000000000000155", x"00003763e74711b0", -80509877, 62);
send(2, x"0000000000000155", x"000033a952a9066c", 161337583, 62);
send(3, x"0000000000000155", x"000030ee9d83d4d0", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ef16807f1", 40296456, 62);
send(1, x"0000000000000155", x"00003763e672c10e", -80509877, 62);
send(2, x"0000000000000155", x"000033a947aa8b6a", 161337583, 62);
send(3, x"0000000000000155", x"000030eea7b9c34a", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ef029ea50", 40296456, 62);
send(1, x"0000000000000155", x"00003763e59e7c65", -80509877, 62);
send(2, x"0000000000000155", x"000033a93cac1367", 161337583, 62);
send(3, x"0000000000000155", x"000030eeb1efbdbe", 120539330, 62);
send(0, x"0000000000000155", x"00002d0eeeebd5aa", 40296456, 62);
send(1, x"0000000000000155", x"00003763e4ca43b6", -80509877, 62);
send(2, x"0000000000000155", x"000033a931ada161", 161337583, 62);
send(3, x"0000000000000155", x"000030eebc25c12e", 120539330, 62);
send(0, x"0000000000000155", x"00002d0eedadcffc", 40296456, 62);
send(1, x"0000000000000155", x"00003763e3f61cff", -80509877, 62);
send(2, x"0000000000000155", x"000033a926af3856", 161337583, 62);
send(3, x"0000000000000155", x"000030eec65bcd99", 120539330, 62);
send(0, x"0000000000000155", x"00002d0eec6fd04c", 40296456, 62);
send(1, x"0000000000000155", x"00003763e3220540", -80509877, 62);
send(2, x"0000000000000155", x"000033a91bb0d549", 161337583, 62);
send(3, x"0000000000000155", x"000030eed091e2ff", 120539330, 62);
send(0, x"0000000000000255", x"00002d0eeb31df94", 40296456, 62);
send(1, x"0000000000000255", x"00003763e24dfc79", -80509877, 62);
send(2, x"0000000000000255", x"000033a910b27b37", 161337583, 62);
send(3, x"0000000000000255", x"000030eedac8075e", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ee9f3f4d9", 40296456, 62);
send(1, x"0000000000000155", x"00003763e179ffad", -80509877, 62);
send(2, x"0000000000000155", x"000033a905b42125", 161337583, 62);
send(3, x"0000000000000155", x"000030eee4fe31ba", 120539330, 62);
send(0, x"000000000000031f", x"00002d0ee8b61916", 40296456, 62);
send(1, x"000000000000031f", x"00003763e0a614d7", -80509877, 62);
send(2, x"000000000000031f", x"000033a8fab5d00e", 161337583, 62);
send(3, x"000000000000031f", x"000030eeef346512", 120539330, 62);
send(0, x"00000000000000ae", x"00002d0ee778494e", 40296456, 62);
send(1, x"00000000000000ae", x"00003763dfd235fc", -80509949, 62);
send(2, x"00000000000000ae", x"000033a8efb784f5", 161337583, 62);
send(3, x"00000000000000ae", x"000030eef96aa164", 120539330, 62);
send(0, x"00000000000001a4", x"00002d0ee63a8281", 40296456, 62);
send(1, x"00000000000001a4", x"00003763defe631b", -80509949, 62);
send(2, x"00000000000001a4", x"000033a8e4b93fd8", 161337583, 62);
send(3, x"00000000000001a4", x"000030ef03a0e9b2", 120539330, 62);
send(0, x"0000000000000196", x"00002d0ee4fcc7ae", 40296456, 62);
send(1, x"0000000000000196", x"00003763de2aa52f", -80509949, 62);
send(2, x"0000000000000196", x"000033a8d9bb00b9", 161337583, 62);
send(3, x"0000000000000196", x"000030ef0dd73afa", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ee3bf15d6", 40296456, 62);
send(1, x"0000000000000155", x"00003763dd56f33d", -80509949, 62);
send(2, x"0000000000000155", x"000033a8cebcc797", 161337583, 62);
send(3, x"0000000000000155", x"000030ef180d953e", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ee2816ff9", 40296456, 62);
send(1, x"0000000000000155", x"00003763dc834d45", -80509949, 62);
send(2, x"0000000000000155", x"000033a8c3be9471", 161337583, 62);
send(3, x"0000000000000155", x"000030ef2243f87e", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ee143d615", 40296456, 62);
send(1, x"0000000000000155", x"00003763dbafb645", -80509949, 62);
send(2, x"0000000000000155", x"000033a8b8c06749", 161337583, 62);
send(3, x"0000000000000155", x"000030ef2c7a67b7", 120539330, 62);
send(0, x"0000000000000155", x"00002d0ee006482b", 40296456, 62);
send(1, x"0000000000000155", x"00003763dadc313d", -80509949, 62);
send(2, x"0000000000000155", x"000033a8adc2431b", 161337511, 62);
send(3, x"0000000000000155", x"000030ef36b0dfec", 120539330, 62);
send(0, x"0000000000000155", x"00002d0edec8c33e", 40296456, 62);
send(1, x"0000000000000155", x"00003763da08bb2d", -80509949, 62);
send(2, x"0000000000000155", x"000033a8a2c421ed", 161337511, 62);
send(3, x"0000000000000155", x"000030ef40e7641b", 120539330, 62);
send(0, x"0000000000000155", x"00002d0edd8b474b", 40296385, 62);
send(1, x"0000000000000155", x"00003763d9354e18", -80509949, 62);
send(2, x"0000000000000155", x"000033a897c606bc", 161337511, 62);
send(3, x"0000000000000155", x"000030ef4b1dee47", 120539330, 62);
send(0, x"0000000000000155", x"00002d0edc4dd753", 40296385, 62);
send(1, x"0000000000000155", x"00003763d861f5f9", -80509949, 62);
send(2, x"0000000000000155", x"000033a88cc7f485", 161337511, 62);
send(3, x"0000000000000155", x"000030ef5554816e", 120539259, 62);
send(0, x"0000000000000155", x"00002d0edb107653", 40296385, 62);
send(1, x"0000000000000155", x"00003763d78ea9d4", -80509949, 62);
send(2, x"0000000000000155", x"000033a881c9e84d", 161337511, 62);
send(3, x"0000000000000155", x"000030ef5f8b2090", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ed9d31b50", 40296385, 62);
send(1, x"0000000000000155", x"00003763d6bb69a9", -80509949, 62);
send(2, x"0000000000000155", x"000033a876cbdf12", 161337511, 62);
send(3, x"0000000000000155", x"000030ef69c1c8ad", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ed895cf45", 40296385, 62);
send(1, x"0000000000000155", x"00003763d5e83b75", -80509949, 62);
send(2, x"0000000000000155", x"000033a86bcddbd4", 161337511, 62);
send(3, x"0000000000000155", x"000030ef73f87cc4", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ed7588c36", 40296385, 62);
send(1, x"0000000000000155", x"00003763d5151c3a", -80510020, 62);
send(2, x"0000000000000155", x"000033a860cfe192", 161337511, 62);
send(3, x"0000000000000155", x"000030ef7e2f36d8", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ed61b5521", 40296385, 62);
send(1, x"0000000000000155", x"00003763d44208f8", -80510020, 62);
send(2, x"0000000000000155", x"000033a855d1ea4f", 161337511, 62);
send(3, x"0000000000000155", x"000030ef8865fce6", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ed4de2707", 40296385, 62);
send(1, x"0000000000000155", x"00003763d36f04af", -80510020, 62);
send(2, x"0000000000000155", x"000033a84ad3ff06", 161337511, 62);
send(3, x"0000000000000155", x"000030ef929ccbf0", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ed3a107e7", 40296385, 62);
send(1, x"0000000000000155", x"00003763d29c125d", -80510020, 62);
send(2, x"0000000000000155", x"000033a83fd616bb", 161337511, 62);
send(3, x"0000000000000155", x"000030ef9cd3a3f5", 120539259, 62);
send(0, x"00000000000002a5", x"00002d0ed263eec3", 40296385, 62);
send(1, x"00000000000002a5", x"00003763d1c92c05", -80510020, 62);
send(2, x"00000000000002a5", x"000033a834d8346c", 161337511, 62);
send(3, x"00000000000002a5", x"000030efa70a8af2", 120539259, 62);
send(0, x"00000000000002aa", x"00002d0ed126e198", 40296385, 62);
send(1, x"00000000000002aa", x"00003763d0f651a7", -80510020, 62);
send(2, x"00000000000002aa", x"000033a829da551d", 161337511, 62);
send(3, x"00000000000002aa", x"000030efb14177ed", 120539259, 62);
send(0, x"000000000000031f", x"00002d0ecfe9e068", 40296385, 62);
send(1, x"000000000000031f", x"00003763d0238940", -80510020, 62);
send(2, x"000000000000031f", x"000033a81edc7ec9", 161337511, 62);
send(3, x"000000000000031f", x"000030efbb786de3", 120539259, 62);
send(0, x"00000000000000ae", x"00002d0eceaceb33", 40296385, 62);
send(1, x"00000000000000ae", x"00003763cf50cfd1", -80510020, 62);
send(2, x"00000000000000ae", x"000033a813deb171", 161337511, 62);
send(3, x"00000000000000ae", x"000030efc5af6cd4", 120539259, 62);
send(0, x"00000000000001a4", x"00002d0ecd6ffef8", 40296385, 62);
send(1, x"00000000000001a4", x"00003763ce7e225d", -80510020, 62);
send(2, x"00000000000001a4", x"000033a808e0e418", 161337511, 62);
send(3, x"00000000000001a4", x"000030efcfe677c0", 120539259, 62);
send(0, x"00000000000002a6", x"00002d0ecc331eb8", 40296385, 62);
send(1, x"00000000000002a6", x"00003763cdab86e0", -80510020, 62);
send(2, x"00000000000002a6", x"000033a7fde322ba", 161337511, 62);
send(3, x"00000000000002a6", x"000030efda1d88a8", 120539259, 62);
send(0, x"00000000000002aa", x"00002d0ecaf64a71", 40296385, 62);
send(1, x"00000000000002aa", x"00003763ccd8fa5a", -80510020, 62);
send(2, x"00000000000002aa", x"000033a7f2e5645a", 161337511, 62);
send(3, x"00000000000002aa", x"000030efe454a58b", 120539259, 62);
send(0, x"0000000000000169", x"00002d0ec9b98225", 40296385, 62);
send(1, x"0000000000000169", x"00003763cc0676d1", -80510020, 62);
send(2, x"0000000000000169", x"000033a7e7e7abf7", 161337511, 62);
send(3, x"0000000000000169", x"000030efee8bce67", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ec87cc2d4", 40296313, 62);
send(1, x"0000000000000155", x"00003763cb34053f", -80510020, 62);
send(2, x"0000000000000155", x"000033a7dce9f991", 161337511, 62);
send(3, x"0000000000000155", x"000030eff8c2fd41", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ec7400f7c", 40296313, 62);
send(1, x"0000000000000155", x"00003763ca61a5a3", -80510092, 62);
send(2, x"0000000000000155", x"000033a7d1ec5026", 161337511, 62);
send(3, x"0000000000000155", x"000030f002fa3814", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ec6036521", 40296313, 62);
send(1, x"0000000000000155", x"00003763c98f5202", -80510092, 62);
send(2, x"0000000000000155", x"000033a7c6eeacb9", 161337511, 62);
send(3, x"0000000000000155", x"000030f00d317ee1", 120539259, 62);
send(0, x"0000000000000155", x"00002d0ec4c6c3c1", 40296313, 62);
send(1, x"0000000000000155", x"00003763c8bd0a5a", -80510092, 62);
send(2, x"0000000000000155", x"000033a7bbf1094b", 161337511, 62);
send(3, x"0000000000000155", x"000030f01768cbac", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ec38a315a", 40296313, 62);
send(1, x"0000000000000155", x"00003763c7ead4a9", -80510092, 62);
send(2, x"0000000000000155", x"000033a7b0f371d8", 161337511, 62);
send(3, x"0000000000000155", x"000030f021a02172", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ec24daaec", 40296313, 62);
send(1, x"0000000000000155", x"00003763c718aaf3", -80510092, 62);
send(2, x"0000000000000155", x"000033a7a5f5e061", 161337511, 62);
send(3, x"0000000000000155", x"000030f02bd78332", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ec1112d7a", 40296313, 62);
send(1, x"0000000000000155", x"00003763c6469035", -80510092, 62);
send(2, x"0000000000000155", x"000033a79af851e9", 161337511, 62);
send(3, x"0000000000000155", x"000030f0360eedee", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ebfd4b903", 40296313, 62);
send(1, x"0000000000000155", x"00003763c574876e", -80510092, 62);
send(2, x"0000000000000155", x"000033a78ffacc6d", 161337511, 62);
send(3, x"0000000000000155", x"000030f0404661a5", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ebe985386", 40296313, 62);
send(1, x"0000000000000155", x"00003763c4a28aa1", -80510092, 62);
send(2, x"0000000000000155", x"000033a784fd4ced", 161337511, 62);
send(3, x"0000000000000155", x"000030f04a7de156", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ebd5bf703", 40296313, 62);
send(1, x"0000000000000155", x"00003763c3d099ce", -80510092, 62);
send(2, x"0000000000000155", x"000033a779ffd06c", 161337511, 62);
send(3, x"0000000000000155", x"000030f054b56a02", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ebc1fa67a", 40296313, 62);
send(1, x"0000000000000155", x"00003763c2febaf2", -80510092, 62);
send(2, x"0000000000000155", x"000033a76f025ce7", 161337511, 62);
send(3, x"0000000000000155", x"000030f05eecfbaa", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ebae35eed", 40296313, 62);
send(1, x"0000000000000155", x"00003763c22ceb0e", -80510092, 62);
send(2, x"0000000000000155", x"000033a76404f25d", 161337439, 62);
send(3, x"0000000000000155", x"000030f06924964d", 120539187, 62);
send(0, x"0000000000000195", x"00002d0eb9a7235b", 40296313, 62);
send(1, x"0000000000000195", x"00003763c15b2a24", -80510092, 62);
send(2, x"0000000000000195", x"000033a759078ad1", 161337439, 62);
send(3, x"0000000000000195", x"000030f0735c3ceb", 120539187, 62);
send(0, x"00000000000002aa", x"00002d0eb86af0c3", 40296313, 62);
send(1, x"00000000000002aa", x"00003763c0897532", -80510092, 62);
send(2, x"00000000000002aa", x"000033a74e0a2644", 161337439, 62);
send(3, x"00000000000002aa", x"000030f07d93ec84", 120539187, 62);
send(0, x"000000000000031f", x"00002d0eb72eca25", 40296313, 62);
send(1, x"000000000000031f", x"00003763bfb7d239", -80510164, 62);
send(2, x"000000000000031f", x"000033a7430ccdb1", 161337439, 62);
send(3, x"000000000000031f", x"000030f087cba519", 120539187, 62);
send(0, x"00000000000000ae", x"00002d0eb5f2af82", 40296313, 62);
send(1, x"00000000000000ae", x"00003763bee63b39", -80510164, 62);
send(2, x"00000000000000ae", x"000033a7380f781d", 161337439, 62);
send(3, x"00000000000000ae", x"000030f0920366a8", 120539187, 62);
send(0, x"00000000000001a4", x"00002d0eb4b6a0d9", 40296313, 62);
send(1, x"00000000000001a4", x"00003763be14b331", -80510164, 62);
send(2, x"00000000000001a4", x"000033a72d122885", 161337439, 62);
send(3, x"00000000000001a4", x"000030f09c3b3134", 120539187, 62);
send(0, x"00000000000001a6", x"00002d0eb37a9e29", 40296242, 62);
send(1, x"00000000000001a6", x"00003763bd433a22", -80510164, 62);
send(2, x"00000000000001a6", x"000033a72214deeb", 161337439, 62);
send(3, x"00000000000001a6", x"000030f0a67307ba", 120539187, 62);
send(0, x"0000000000000155", x"00002d0eb23ea475", 40296242, 62);
send(1, x"0000000000000155", x"00003763bc71d00c", -80510164, 62);
send(2, x"0000000000000155", x"000033a717179e4c", 161337439, 62);
send(3, x"0000000000000155", x"000030f0b0aae73b", 120539187, 62);
send(0, x"0000000000000155", x"00002d0eb102b3bd", 40296242, 62);
send(1, x"0000000000000155", x"00003763bba071ef", -80510164, 62);
send(2, x"0000000000000155", x"000033a70c1a60ab", 161337439, 62);
send(3, x"0000000000000155", x"000030f0bae2cfb7", 120539187, 62);
send(0, x"0000000000000155", x"00002d0eafc6d1fd", 40296242, 62);
send(1, x"0000000000000155", x"00003763bacf25ca", -80510164, 62);
send(2, x"0000000000000155", x"000033a7011d2908", 161337439, 62);
send(3, x"0000000000000155", x"000030f0c51ac12f", 120539187, 62);
send(0, x"0000000000000155", x"00002d0eae8af938", 40296242, 62);
send(1, x"0000000000000155", x"00003763b9fde89c", -80510164, 62);
send(2, x"0000000000000155", x"000033a6f61ffa60", 161337439, 62);
send(3, x"0000000000000155", x"000030f0cf52bea1", 120539187, 62);
send(0, x"0000000000000155", x"00002d0ead4f2c6e", 40296242, 62);
send(1, x"0000000000000155", x"00003763b92cb769", -80510164, 62);
send(2, x"0000000000000155", x"000033a6eb22d1b5", 161337439, 62);
send(3, x"0000000000000155", x"000030f0d98ac80d", 120539116, 62);
send(0, x"0000000000000155", x"00002d0eac1365a0", 40296242, 62);
send(1, x"0000000000000155", x"00003763b85b952f", -80510164, 62);
send(2, x"0000000000000155", x"000033a6e025ac08", 161337439, 62);
send(3, x"0000000000000155", x"000030f0e3c2d776", 120539116, 62);
send(0, x"0000000000000155", x"00002d0eaad7adcb", 40296242, 62);
send(1, x"0000000000000155", x"00003763b78a84ec", -80510164, 62);
send(2, x"0000000000000155", x"000033a6d5288f57", 161337439, 62);
send(3, x"0000000000000155", x"000030f0edfaefda", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea99c01f0", 40296242, 62);
send(1, x"0000000000000155", x"00003763b6b980a2", -80510164, 62);
send(2, x"0000000000000155", x"000033a6ca2b78a3", 161337439, 62);
send(3, x"0000000000000155", x"000030f0f8331439", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea8605f11", 40296242, 62);
send(1, x"0000000000000155", x"00003763b5e88853", -80510235, 62);
send(2, x"0000000000000155", x"000033a6bf2e64ed", 161337439, 62);
send(3, x"0000000000000155", x"000030f1026b4193", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea724c82b", 40296242, 62);
send(1, x"0000000000000155", x"00003763b517a1fa", -80510235, 62);
send(2, x"0000000000000155", x"000033a6b4315a33", 161337439, 62);
send(3, x"0000000000000155", x"000030f10ca377e9", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea5e93d40", 40296242, 62);
send(1, x"0000000000000155", x"00003763b446ca9a", -80510235, 62);
send(2, x"0000000000000155", x"000033a6a9345577", 161337439, 62);
send(3, x"0000000000000155", x"000030f116dbb73a", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea4adbb50", 40296242, 62);
send(1, x"0000000000000155", x"00003763b375ff34", -80510235, 62);
send(2, x"0000000000000155", x"000033a69e3753b8", 161337439, 62);
send(3, x"0000000000000155", x"000030f121140285", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea372455a", 40296242, 62);
send(1, x"0000000000000155", x"00003763b2a545c5", -80510235, 62);
send(2, x"0000000000000155", x"000033a6933a5df4", 161337439, 62);
send(3, x"0000000000000155", x"000030f12b4c56cb", 120539116, 62);
send(0, x"0000000000000155", x"00002d0ea236db5e", 40296242, 62);
send(1, x"0000000000000155", x"00003763b1d49850", -80510235, 62);
send(2, x"0000000000000155", x"000033a6883d6b2d", 161337439, 62);
send(3, x"0000000000000155", x"000030f13584b40d", 120539116, 62);
send(0, x"0000000000000295", x"00002d0ea0fb7a5d", 40296242, 62);
send(1, x"0000000000000295", x"00003763b103f9d4", -80510235, 62);
send(2, x"0000000000000295", x"000033a67d408163", 161337439, 62);
send(3, x"0000000000000295", x"000030f13fbd1d49", 120539116, 62);
send(0, x"00000000000002aa", x"00002d0e9fc02258", 40296242, 62);
send(1, x"00000000000002aa", x"00003763b0336a50", -80510235, 62);
send(2, x"00000000000002aa", x"000033a672439799", 161337439, 62);
send(3, x"00000000000002aa", x"000030f149f58c82", 120539116, 62);
send(0, x"000000000000031f", x"00002d0e9e84d94c", 40296170, 62);
send(1, x"000000000000031f", x"00003763af62e9c4", -80510235, 62);
send(2, x"000000000000031f", x"000033a66746b9c8", 161337439, 62);
send(3, x"000000000000031f", x"000030f1542e07b5", 120539116, 62);
send(0, x"00000000000000ae", x"00002d0e9d49993a", 40296170, 62);
send(1, x"00000000000000ae", x"00003763ae927831", -80510235, 62);
send(2, x"00000000000000ae", x"000033a65c49def6", 161337439, 62);
send(3, x"00000000000000ae", x"000030f15e668be4", 120539116, 62);
send(0, x"00000000000001a4", x"00002d0e9c0e6524", 40296170, 62);
send(1, x"00000000000001a4", x"00003763adc21298", -80510235, 62);
send(2, x"00000000000001a4", x"000033a6514d0a21", 161337439, 62);
send(3, x"00000000000001a4", x"000030f1689f190d", 120539116, 62);
send(0, x"0000000000000166", x"00002d0e9ad33d07", 40296170, 62);
send(1, x"0000000000000166", x"00003763acf1bef6", -80510235, 62);
send(2, x"0000000000000166", x"000033a646503e48", 161337439, 62);
send(3, x"0000000000000166", x"000030f172d7b232", 120539116, 62);
send(0, x"0000000000000155", x"00002d0e99981de5", 40296170, 62);
send(1, x"0000000000000155", x"00003763ac217a4d", -80510235, 62);
send(2, x"0000000000000155", x"000033a63b53756c", 161337439, 62);
send(3, x"0000000000000155", x"000030f17d105451", 120539116, 62);
send(0, x"0000000000000165", x"00002d0e985d0abe", 40296170, 62);
send(1, x"0000000000000165", x"00003763ab513e9f", -80510307, 62);
send(2, x"0000000000000165", x"000033a63056b28f", 161337439, 62);
send(3, x"0000000000000165", x"000030f18748ff6c", 120539116, 62);
send(0, x"0000000000000155", x"00002d0e97220390", 40296170, 62);
send(1, x"0000000000000155", x"00003763aa8117e6", -80510307, 62);
send(2, x"0000000000000155", x"000033a62559f8ac", 161337439, 62);
send(3, x"0000000000000155", x"000030f19181b383", 120539116, 62);
send(0, x"0000000000000155", x"00002d0e95e7055e", 40296170, 62);
send(1, x"0000000000000155", x"00003763a9b0fd28", -80510307, 62);
send(2, x"0000000000000155", x"000033a61a5d44c7", 161337368, 62);
send(3, x"0000000000000155", x"000030f19bba7095", 120539116, 62);
send(0, x"0000000000000155", x"00002d0e94ac1326", 40296170, 62);
send(1, x"0000000000000155", x"00003763a8e0f161", -80510307, 62);
send(2, x"0000000000000155", x"000033a60f6096de", 161337368, 62);
send(3, x"0000000000000155", x"000030f1a5f33c9f", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e937129ea", 40296170, 62);
send(1, x"0000000000000155", x"00003763a810f196", -80510307, 62);
send(2, x"0000000000000155", x"000033a60463ebf4", 161337368, 62);
send(3, x"0000000000000155", x"000030f1b02c0ea6", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e92364ca7", 40296170, 62);
send(1, x"0000000000000155", x"00003763a74103c1", -80510307, 62);
send(2, x"0000000000000155", x"000033a5f9674a06", 161337368, 62);
send(3, x"0000000000000155", x"000030f1ba64e9aa", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e90fb7b5e", 40296170, 62);
send(1, x"0000000000000155", x"00003763a67124e4", -80510307, 62);
send(2, x"0000000000000155", x"000033a5ee6aae14", 161337368, 62);
send(3, x"0000000000000155", x"000030f1c49dd0a6", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e8fc0b610", 40296170, 62);
send(1, x"0000000000000155", x"00003763a5a15202", -80510307, 62);
send(2, x"0000000000000155", x"000033a5e36e1820", 161337368, 62);
send(3, x"0000000000000155", x"000030f1ced6bda1", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e8e85f9bd", 40296170, 62);
send(1, x"0000000000000155", x"00003763a4d19116", -80510307, 62);
send(2, x"0000000000000155", x"000033a5d8718828", 161337368, 62);
send(3, x"0000000000000155", x"000030f1d90fb695", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e8d4b4964", 40296170, 62);
send(1, x"0000000000000155", x"00003763a401dc24", -80510307, 62);
send(2, x"0000000000000155", x"000033a5cd74fe2e", 161337368, 62);
send(3, x"0000000000000155", x"000030f1e348bb82", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e8c10a505", 40296170, 62);
send(1, x"0000000000000155", x"00003763a332332d", -80510307, 62);
send(2, x"0000000000000155", x"000033a5c2787a30", 161337368, 62);
send(3, x"0000000000000155", x"000030f1ed81c66d", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e8ad609a2", 40296170, 62);
send(1, x"0000000000000155", x"00003763a2629f2b", -80510307, 62);
send(2, x"0000000000000155", x"000033a5b77bfc30", 161337368, 62);
send(3, x"0000000000000155", x"000030f1f7badd53", 120539044, 62);
send(0, x"0000000000000155", x"00002d0e899b7a38", 40296098, 62);
send(1, x"0000000000000155", x"00003763a1931723", -80510307, 62);
send(2, x"0000000000000155", x"000033a5ac7f872a", 161337368, 62);
send(3, x"0000000000000155", x"000030f201f3fd33", 120539044, 62);
send(0, x"0000000000000255", x"00002d0e8860f6c9", 40296098, 62);
send(1, x"0000000000000255", x"00003763a0c39e14", -80510378, 62);
send(2, x"0000000000000255", x"000033a5a1831524", 161337368, 62);
send(3, x"0000000000000255", x"000030f20c2d290e", 120539044, 62);
send(0, x"00000000000002aa", x"00002d0e87267956", 40296098, 62);
send(1, x"00000000000002aa", x"000037639ff430fe", -80510378, 62);
send(2, x"00000000000002aa", x"000033a59686a91b", 161337368, 62);
send(3, x"00000000000002aa", x"000030f216665ae5", 120539044, 62);
send(0, x"000000000000031f", x"00002d0e85ec0adc", 40296098, 62);
send(1, x"000000000000031f", x"000037639f24d2e1", -80510378, 62);
send(2, x"000000000000031f", x"000033a58b8a460d", 161337368, 62);
send(3, x"000000000000031f", x"000030f2209f98b7", 120539044, 62);
send(0, x"00000000000000ae", x"00002d0e84b1a55e", 40296098, 62);
send(1, x"00000000000000ae", x"000037639e5586bb", -80510378, 62);
send(2, x"00000000000000ae", x"000033a5808de8fc", 161337368, 62);
send(3, x"00000000000000ae", x"000030f22ad8dc85", 120539044, 62);
send(0, x"00000000000001a4", x"00002d0e83774ed8", 40296098, 62);
send(1, x"00000000000001a4", x"000037639d86468f", -80510378, 62);
send(2, x"00000000000001a4", x"000033a575918ee9", 161337368, 62);
send(3, x"00000000000001a4", x"000030f235122f4c", 120539044, 62);
send(0, x"0000000000000266", x"00002d0e823d014d", 40296098, 62);
send(1, x"0000000000000266", x"000037639cb7155c", -80510378, 62);
send(2, x"0000000000000266", x"000033a56a953ad4", 161337368, 62);
send(3, x"0000000000000266", x"000030f23f4b8810", 120539044, 62);
send(0, x"00000000000002aa", x"00002d0e8102bcbe", 40296098, 62);
send(1, x"00000000000002aa", x"000037639be7f321", -80510378, 62);
send(2, x"00000000000002aa", x"000033a55f98efb9", 161337368, 62);
send(3, x"00000000000002aa", x"000030f24984e9cf", 120539044, 62);
send(0, x"00000000000002aa", x"00002d0e7fc88429", 40296098, 62);
send(1, x"00000000000002aa", x"000037639b18dcdf", -80510378, 62);
send(2, x"00000000000002aa", x"000033a5549ca79e", 161337368, 62);
send(3, x"00000000000002aa", x"000030f253be5789", 120539044, 62);
send(0, x"00000000000002aa", x"00002d0e7e8e578e", 40296098, 62);
send(1, x"00000000000002aa", x"000037639a49d896", -80510378, 62);
send(2, x"00000000000002aa", x"000033a549a06b7d", 161337368, 62);
send(3, x"00000000000002aa", x"000030f25df7ce3e", 120539044, 62);
send(0, x"00000000000002aa", x"00002d0e7d5436ed", 40296098, 62);
send(1, x"00000000000002aa", x"00003763997ae344", -80510378, 62);
send(2, x"00000000000002aa", x"000033a53ea4325a", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2683150ed", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e7c1a1f48", 40296098, 62);
send(1, x"00000000000002aa", x"0000376398abfceb", -80510378, 62);
send(2, x"00000000000002aa", x"000033a533a7ff34", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2726adc98", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e7ae0109e", 40296098, 62);
send(1, x"00000000000002aa", x"0000376397dd228c", -80510378, 62);
send(2, x"00000000000002aa", x"000033a528abcf0c", 161337368, 62);
send(3, x"00000000000002aa", x"000030f27ca4713d", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e79a610ec", 40296098, 62);
send(1, x"00000000000002aa", x"00003763970e5726", -80510378, 62);
send(2, x"00000000000002aa", x"000033a51dafaade", 161337368, 62);
send(3, x"00000000000002aa", x"000030f286de0edf", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e786c1a36", 40296098, 62);
send(1, x"00000000000002aa", x"00003763963f9db6", -80510450, 62);
send(2, x"00000000000002aa", x"000033a512b389b0", 161337368, 62);
send(3, x"00000000000002aa", x"000030f29117b57c", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e77322f7a", 40296098, 62);
send(1, x"00000000000002aa", x"000037639570ed42", -80510450, 62);
send(2, x"00000000000002aa", x"000033a507b76b7f", 161337368, 62);
send(3, x"00000000000002aa", x"000030f29b516813", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e75f84db9", 40296098, 62);
send(1, x"00000000000002aa", x"0000376394a24ec5", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4fcbb5948", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2a58b23a6", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e74be77f3", 40296027, 62);
send(1, x"00000000000002aa", x"0000376393d3bf41", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4f1bf4a11", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2afc4e834", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e7384ae26", 40296027, 62);
send(1, x"00000000000002aa", x"0000376393053bb6", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4e6c340d6", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2b9feb5bd", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e724af054", 40296027, 62);
send(1, x"00000000000002aa", x"000037639236ca23", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4dbc74096", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2c4388c42", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e71113b7d", 40296027, 62);
send(1, x"00000000000002aa", x"0000376391686788", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4d0cb4654", 161337368, 62);
send(3, x"00000000000002aa", x"000030f2ce726ec1", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e6fd792a0", 40296027, 62);
send(1, x"00000000000002aa", x"00003763909a10e7", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4c5cf4f10", 161337296, 62);
send(3, x"00000000000002aa", x"000030f2d8ac5d3a", 120538972, 62);
send(0, x"00000000000002aa", x"00002d0e6e9defc0", 40296027, 62);
send(1, x"00000000000002aa", x"000037638fcbc93e", -80510450, 62);
send(2, x"00000000000002aa", x"000033a4bad35dc9", 161337296, 62);
send(3, x"00000000000002aa", x"000030f2e2e651b0", 120538972, 62);
send(0, x"000000000000031f", x"00002d0e6d645ed7", 40296027, 62);
send(1, x"000000000000031f", x"000037638efd908e", -80510450, 62);
send(2, x"000000000000031f", x"000033a4afd7757d", 161337296, 62);
send(3, x"000000000000031f", x"000030f2ed204f21", 120538972, 62);
send(0, x"00000000000000ae", x"00002d0e6c2ad3eb", 40296027, 62);
send(1, x"00000000000000ae", x"000037638e2f66d7", -80510450, 62);
send(2, x"00000000000000ae", x"000033a4a4db932f", 161337296, 62);
send(3, x"00000000000000ae", x"000030f2f75a588d", 120538972, 62);
send(0, x"00000000000001a4", x"00002d0e6af157f8", 40296027, 62);
send(1, x"00000000000001a4", x"000037638d614919", -80510450, 62);
send(2, x"00000000000001a4", x"000033a499dfb3de", 161337296, 62);
send(3, x"00000000000001a4", x"000030f301946af4", 120538972, 62);
send(0, x"00000000000001aa", x"00002d0e69b7e500", 40296027, 62);
send(1, x"00000000000001aa", x"000037638c933d53", -80510450, 62);
send(2, x"00000000000001aa", x"000033a48ee3e089", 161337296, 62);
send(3, x"00000000000001aa", x"000030f30bce8657", 120538972, 62);
send(0, x"0000000000000295", x"00002d0e687e7e02", 40296027, 62);
send(1, x"0000000000000295", x"000037638bc54085", -80510522, 62);
send(2, x"0000000000000295", x"000033a483e81031", 161337296, 62);
send(3, x"0000000000000295", x"000030f31608adb3", 120538972, 62);
send(0, x"000000000000015a", x"00002d0e67451fff", 40296027, 62);
send(1, x"000000000000015a", x"000037638af74fb0", -80510522, 62);
send(2, x"000000000000015a", x"000033a478ec42d8", 161337296, 62);
send(3, x"000000000000015a", x"000030f32042db0c", 120538972, 62);
send(0, x"0000000000000155", x"00002d0e660bcdf7", 40296027, 62);
send(1, x"0000000000000155", x"000037638a296dd5", -80510522, 62);
send(2, x"0000000000000155", x"000033a46df07e7a", 161337296, 62);
send(3, x"0000000000000155", x"000030f32a7d1460", 120538901, 62);
send(0, x"0000000000000256", x"00002d0e64d287e8", 40296027, 62);
send(1, x"0000000000000156", x"00003763895b9df0", -80510522, 62);
send(2, x"000000000000016a", x"000033a462f4c319", 161337296, 62);
send(3, x"00000000000002aa", x"000030f334b756af", 120538901, 62);
send(0, x"0000000000000159", x"00002d0e63994dd4", 40296027, 62);
send(1, x"0000000000000165", x"00003763888dda06", -80510522, 62);
send(2, x"000000000000029a", x"000033a457f90ab5", 161337296, 62);
send(3, x"00000000000001a9", x"000030f33ef1a4f8", 120538901, 62);
send(0, x"0000000000000295", x"00002d0e626019bc", 40296027, 62);
send(1, x"00000000000002a5", x"0000376387c02216", -80510522, 62);
send(2, x"0000000000000269", x"000033a44cfd584f", 161337296, 62);
send(3, x"0000000000000155", x"000030f3492bfc3d", 120538901, 62);
send(0, x"0000000000000256", x"00002d0e6126f49d", 40296027, 62);
send(1, x"0000000000000266", x"0000376386f27c1c", -80510522, 62);
send(2, x"00000000000001a5", x"000033a44201abe5", 161337296, 62);
send(3, x"0000000000000259", x"000030f353665c7d", 120538901, 62);
send(0, x"0000000000000199", x"00002d0e5fedd87a", 40295955, 62);
send(1, x"0000000000000299", x"000037638624e51b", -80510522, 62);
send(2, x"0000000000000269", x"000033a437060877", 161337296, 62);
send(3, x"00000000000001a6", x"000030f35da0c5b8", 120538901, 62);
send(0, x"00000000000001a5", x"00002d0e5eb4c850", 40295955, 62);
send(1, x"00000000000002aa", x"0000376385575a14", -80510522, 62);
send(2, x"000000000000025a", x"000033a42c0a6808", 161337296, 62);
send(3, x"0000000000000295", x"000030f367db37ef", 120538901, 62);
send(0, x"00000000000001a9", x"00002d0e5d7bc421", 40295955, 62);
send(1, x"00000000000002a5", x"000037638489e104", -80510522, 62);
send(2, x"0000000000000155", x"000033a4210ecd95", 161337296, 62);
send(3, x"0000000000000196", x"000030f37215b620", 120538901, 62);
send(0, x"0000000000000259", x"00002d0e5c42c8ec", 40295955, 62);
send(1, x"0000000000000256", x"0000376383bc76ed", -80510522, 62);
send(2, x"00000000000001aa", x"000033a416133c1e", 161337296, 62);
send(3, x"00000000000002a9", x"000030f37c503a4e", 120538901, 62);
send(0, x"0000000000000269", x"00002d0e5b09dcb1", 40295955, 62);
send(1, x"0000000000000155", x"0000376382ef15d1", -80510522, 62);
send(2, x"00000000000001a5", x"000033a40b17ada6", 161337296, 62);
send(3, x"000000000000016a", x"000030f3868acd75", 120538901, 62);
send(0, x"0000000000000166", x"00002d0e59d0f673", 40295955, 62);
send(1, x"0000000000000165", x"000037638221c6ac", -80510593, 62);
send(2, x"000000000000015a", x"000033a4001c2829", 161337296, 62);
send(3, x"000000000000016a", x"000030f390c56698", 120538901, 62);
send(0, x"0000000000000266", x"00002d0e58981f2d", 40295955, 62);
send(1, x"0000000000000159", x"000037638154897d", -80510593, 62);
send(2, x"0000000000000196", x"000033a3f520a8a9", 161337296, 62);
send(3, x"000000000000016a", x"000030f39b0008b7", 120538901, 62);
send(0, x"00000000000002a9", x"00002d0e575f50e2", 40295955, 62);
send(1, x"0000000000000295", x"000037638087584a", -80510593, 62);
send(2, x"00000000000002a5", x"000033a3ea252f26", 161337296, 62);
send(3, x"0000000000000156", x"000030f3a53ab9cf", 120538901, 62);
send(0, x"00000000000002a5", x"00002d0e56268b93", 40295955, 62);
send(1, x"00000000000002a5", x"000037637fba330f", -80510593, 62);
send(2, x"0000000000000159", x"000033a3df29b8a1", 161337296, 62);
send(3, x"00000000000002a9", x"000030f3af7570e3", 120538901, 62);
send(0, x"000000000000031f", x"00002d0e54edd23e", 40295955, 62);
send(1, x"000000000000031f", x"000037637eed1fcd", -80510593, 62);
send(2, x"000000000000031f", x"000033a3d42e4e17", 161337296, 62);
send(3, x"000000000000031f", x"000030f3b9b030f3", 120538901, 62);
send(0, x"00000000000000ae", x"00002d0e53b524e3", 40295955, 62);
send(1, x"00000000000000ae", x"000037637e201883", -80510593, 62);
send(2, x"00000000000000ae", x"000033a3c932e68b", 161337296, 62);
send(3, x"00000000000000ae", x"000030f3c3eafcfd", 120538901, 62);
send(0, x"00000000000001a4", x"00002d0e527c8382", 40295955, 62);
send(1, x"00000000000001a4", x"000037637d532033", -80510593, 62);
send(2, x"00000000000001a4", x"000033a3be3781fd", 161337296, 62);
send(3, x"00000000000001a4", x"000030f3ce25cf04", 120538901, 62);
send(0, x"000000000000016a", x"00002d0e5143eb1d", 40295955, 62);
send(1, x"000000000000016a", x"000037637c8639da", -80510593, 62);
send(2, x"000000000000016a", x"000033a3b33c2969", 161337296, 62);
send(3, x"000000000000016a", x"000030f3d860ad05", 120538901, 62);
send(0, x"0000000000000155", x"00002d0e500b5eb1", 40295955, 62);
send(1, x"0000000000000155", x"000037637bb95f7a", -80510593, 62);
send(2, x"0000000000000155", x"000033a3a840d3d4", 161337296, 62);
send(3, x"0000000000000155", x"000030f3e29b9402", 120538901, 62);
send(0, x"0000000000000195", x"00002d0e4ed2de40", 40295955, 62);
send(1, x"0000000000000195", x"000037637aec9115", -80510593, 62);
send(2, x"0000000000000195", x"000033a39d45843d", 161337296, 62);
send(3, x"0000000000000195", x"000030f3ecd686f8", 120538829, 62);
send(0, x"00000000000002aa", x"00002d0e4d9a66ca", 40295955, 62);
send(1, x"00000000000002aa", x"000037637a1fd7a5", -80510593, 62);
send(2, x"00000000000002aa", x"000033a3924a3aa2", 161337296, 62);
send(3, x"00000000000002aa", x"000030f3f7117fec", 120538829, 62);
send(0, x"00000000000001aa", x"00002d0e4c61fb4e", 40295955, 62);
send(1, x"0000000000000296", x"0000376379532a2f", -80510593, 62);
send(2, x"00000000000001aa", x"000033a3874efa02", 161337296, 62);
send(3, x"00000000000002aa", x"000030f4014c84d9", 120538829, 62);
send(0, x"00000000000001a5", x"00002d0e4b299bcb", 40295884, 62);
send(1, x"0000000000000265", x"00003763788688b2", -80510593, 62);
send(2, x"0000000000000299", x"000033a37c53bf5f", 161337225, 62);
send(3, x"000000000000015a", x"000030f40b8795c1", 120538829, 62);
send(0, x"0000000000000259", x"00002d0e49f14545", 40295884, 62);
send(1, x"0000000000000296", x"0000376377b9f62f", -80510665, 62);
send(2, x"000000000000019a", x"000033a3715884bd", 161337225, 62);
send(3, x"0000000000000156", x"000030f415c2afa4", 120538829, 62);
send(0, x"0000000000000159", x"00002d0e48b8fab9", 40295884, 62);
send(1, x"0000000000000169", x"0000376376ed75a3", -80510665, 62);
send(2, x"0000000000000269", x"000033a3665d5614", 161337225, 62);
send(3, x"0000000000000295", x"000030f41ffdcf84", 120538829, 62);
send(0, x"000000000000016a", x"00002d0e4780b928", 40295884, 62);
send(1, x"00000000000002a5", x"0000376376210110", -80510665, 62);
send(2, x"00000000000001a5", x"000033a35b622d69", 161337225, 62);
send(3, x"00000000000002a6", x"000030f42a38fb5e", 120538829, 62);
send(0, x"000000000000026a", x"00002d0e4648868f", 40295884, 62);
send(1, x"0000000000000255", x"0000376375549b76", -80510665, 62);
send(2, x"00000000000001aa", x"000033a3506707bc", 161337225, 62);
send(3, x"00000000000002a5", x"000030f434743033", 120538829, 62);
send(0, x"0000000000000295", x"00002d0e45105cf2", 40295884, 62);
send(1, x"000000000000029a", x"00003763748844d4", -80510665, 62);
send(2, x"000000000000025a", x"000033a3456beb0b", 161337225, 62);
send(3, x"000000000000015a", x"000030f43eaf6e04", 120538829, 62);
send(0, x"00000000000002aa", x"00002d0e43d83c51", 40295884, 62);
send(1, x"00000000000001a6", x"0000376373bbfd2c", -80510665, 62);
send(2, x"0000000000000159", x"000033a33a70d456", 161337225, 62);
send(3, x"000000000000026a", x"000030f448eab7cf", 120538829, 62);
send(0, x"00000000000002a5", x"00002d0e42a027a9", 40295884, 62);
send(1, x"000000000000025a", x"0000376372efc47b", -80510665, 62);
send(2, x"000000000000016a", x"000033a32f75c39e", 161337225, 62);
send(3, x"0000000000000166", x"000030f453260a95", 120538829, 62);
send(0, x"0000000000000256", x"00002d0e41681efc", 40295884, 62);
send(1, x"0000000000000296", x"00003763722397c5", -80510665, 62);
send(2, x"0000000000000165", x"000033a3247ab8e4", 161337225, 62);
send(3, x"000000000000029a", x"000030f45d616658", 120538829, 62);
send(0, x"0000000000000265", x"00002d0e40302248", 40295884, 62);
send(1, x"0000000000000199", x"0000376371577d05", -80510665, 62);
send(2, x"0000000000000295", x"000033a3197fb426", 161337225, 62);
send(3, x"0000000000000259", x"000030f4679ccb15", 120538829, 62);
send(0, x"000000000000016a", x"00002d0e3ef82e90", 40295884, 62);
send(1, x"0000000000000156", x"00003763708b713e", -80510665, 62);
send(2, x"0000000000000269", x"000033a30e84b566", 161337225, 62);
send(3, x"0000000000000256", x"000030f471d83bcd", 120538829, 62);
send(0, x"00000000000002a5", x"00002d0e3dc043d4", 40295884, 62);
send(1, x"000000000000029a", x"000037636fbf7171", -80510665, 62);
send(2, x"000000000000016a", x"000033a30389bca3", 161337225, 62);
send(3, x"0000000000000155", x"000030f47c13b580", 120538829, 62);
send(0, x"000000000000031f", x"00002d0e3c886810", 40295884, 62);
send(1, x"000000000000031f", x"000037636ef3809d", -80510665, 62);
send(2, x"000000000000031f", x"000033a2f88ec9dc", 161337225, 62);
send(3, x"000000000000031f", x"000030f4864f382e", 120538829, 62);
send(0, x"00000000000000ae", x"00002d0e3b509547", 40295884, 62);
send(1, x"00000000000000ae", x"000037636e279ec0", -80510665, 62);
send(2, x"00000000000000ae", x"000033a2ed93e011", 161337225, 62);
send(3, x"00000000000000ae", x"000030f4908ac3d8", 120538829, 62);
send(0, x"00000000000001a4", x"00002d0e3a18ce79", 40295884, 62);
send(1, x"00000000000001a4", x"000037636d5bcbdd", -80510736, 62);
send(2, x"00000000000001a4", x"000033a2e298f944", 161337225, 62);
send(3, x"00000000000001a4", x"000030f49ac65b7c", 120538829, 62);
send(0, x"000000000000026a", x"00002d0e38e113a4", 40295884, 62);
send(1, x"000000000000026a", x"000037636c9007f2", -80510736, 62);
send(2, x"000000000000026a", x"000033a2d79e1875", 161337225, 62);
send(3, x"000000000000026a", x"000030f4a501f91d", 120538829, 62);
send(0, x"0000000000000155", x"00002d0e37a961cb", 40295884, 62);
send(1, x"0000000000000155", x"000037636bc45300", -80510736, 62);
send(2, x"0000000000000155", x"000033a2cca340a1", 161337225, 62);
send(3, x"00000000000002a9", x"000030f4af3da2b8", 120538829, 62);
send(0, x"0000000000000155", x"00002d0e3671bbec", 40295812, 62);
send(1, x"0000000000000155", x"000037636af8aa07", -80510736, 62);
send(2, x"0000000000000155", x"000033a2c1a86bcb", 161337225, 62);
send(3, x"00000000000002aa", x"000030f4b979554f", 120538758, 62);
send(0, x"00000000000002a9", x"00002d0e353a2207", 40295812, 62);
send(1, x"0000000000000156", x"000037636a2d1007", -80510736, 62);
send(2, x"0000000000000156", x"000033a2b6ad9ff1", 161337225, 62);
send(3, x"0000000000000156", x"000030f4c3b513df", 120538758, 62);
send(0, x"000000000000016a", x"00002d0e3402911e", 40295812, 62);
send(1, x"0000000000000255", x"00003763696187fe", -80510736, 62);
send(2, x"0000000000000155", x"000033a2abb2da15", 161337225, 62);
send(3, x"0000000000000269", x"000030f4cdf0d86d", 120538758, 62);
send(0, x"00000000000001aa", x"00002d0e32cb0c2e", 40295812, 62);
send(1, x"0000000000000165", x"0000376368960bef", -80510736, 62);
send(2, x"00000000000002a6", x"000033a2a0b81a35", 161337225, 62);
send(3, x"0000000000000155", x"000030f4d82cabf3", 120538758, 62);
send(0, x"00000000000001aa", x"00002d0e3193903a", 40295812, 62);
send(1, x"0000000000000199", x"0000376367ca9ed9", -80510736, 62);
send(2, x"0000000000000199", x"000033a295bd5d53", 161337225, 62);
send(3, x"0000000000000295", x"000030f4e2688576", 120538758, 62);
send(0, x"0000000000000166", x"00002d0e305c2040", 40295812, 62);
send(1, x"0000000000000165", x"0000376366ff40ba", -80510736, 62);
send(2, x"0000000000000196", x"000033a28ac2a96d", 161337225, 62);
send(3, x"00000000000002a9", x"000030f4eca46af3", 120538758, 62);
send(0, x"0000000000000266", x"00002d0e2f24bc40", 40295812, 62);
send(1, x"0000000000000195", x"000037636633f195", -80510736, 62);
send(2, x"0000000000000199", x"000033a27fc7fb84", 161337225, 62);
send(3, x"0000000000000295", x"000030f4f6e0566d", 120538758, 62);
        
      loop
        word <= (others => '0');
        wait until rising_edge(send_done);
        word <= (others => '1');
        wait until rising_edge(send_done);
      end loop;
      
    end process;

end;
