library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package input is
  
  constant inputFrameSatCount : integer := 1;
  
  type inputTable is array(0 to 100 - 1) of std_logic_vector(176-1 downto 0);
  constant inputSeq : inputTable := (
    x"0004000000000000b41a0000000000000000000000ff",
    x"00040000000001e90fc30000000000000000000000ff",
    x"000400000000017e1f9f0000000000000000000000ff",
    x"00040000000000d604000000000000000000000000ff",
    x"00040000000000df7fff0000000000000000000000ff",
    x"000400000000000802630000000000000000000000ff",
    x"00040000000000fffbe10000000000000000000000ff",
    x"000400000000000afc9f0000000000000000000000ff",
    x"000400000000014a68100000000000000000000000ff",
    x"000400000000007c7bff0000000000000000000000ff",
    x"00040000000001dc901a0000000000000000000000ff",
    x"000400000000013596980000000000000000000000ff",
    x"00040000000001a475f30000000000000000000000ff",
    x"000400000000014542e80000000000000000000000ff",
    x"0004000000000193e4950000000000000000000000ff",
    x"000400000000004f78430000000000000000000000ff",
    x"00040000000000880dcc0000000000000000000000ff",
    x"000400000000007701f30000000000000000000000ff",
    x"000400000000009b1c060000000000000000000000ff",
    x"00040000000000092e0a0000000000000000000000ff",
    x"00040000000000001c1a0000000000000000000000ff",
    x"00040000000001fc20c30000000000000000000000ff",
    x"00040000000000152f9f0000000000000000000000ff",
    x"000400000000010604000000000000000000000000ff",
    x"000400000000003f7ffd0000000000000000000000ff",
    x"000400000000000800dc0000000000000000000000ff",
    x"00040000000000ffcea60000000000000000000000ff",
    x"000400000000000448ff0000000000000000000000ff",
    x"000400000000012b2c100000000000000000000000ff",
    x"00040000000000717bff0000000000000000000000ff",
    x"0004000000000002e01a0000000000000000000000ff",
    x"00040000000001e180000000000000000000000000ff",
    x"00040000000001afffff0000000000000000000000ff",
    x"000400000000000000070000000000000000000000ff",
    x"00040000000001ffff410000000000000000000000ff",
    x"0004000000000000071f0000000000000000000000ff",
    x"00040000000001fe14000000000000000000000000ff",
    x"000400000000003f7fff0000000000000000000000ff",
    x"000400000000003000000000000000000000000000ff",
    x"00040000000001fffffe0000000000000000000000ff",
    x"0004000000000000041a0000000000000000000000ff",
    x"00040000000001ff1b030000000000000000000000ff",
    x"000400000000001d379f0000000000000000000000ff",
    x"00040000000000f504000000000000000000000000ff",
    x"000400000000003f7ffd0000000000000000000000ff",
    x"000400000000000800660000000000000000000000ff",
    x"00040000000000fff37e0000000000000000000000ff",
    x"0004000000000000f5ff0000000000000000000000ff",
    x"00040000000001e86c100000000000000000000000ff",
    x"000400000000002c7bff0000000000000000000000ff",
    x"0004000000000000101a0000000000000000000000ff",
    x"00040000000001fd8c000000000000000000000000ff",
    x"0004000000000040ffff0000000000000000000000ff",
    x"00040000000001b000000000000000000000000000ff",
    x"00040000000001fffff70000000000000000000000ff",
    x"000400000000000001820000000000000000000000ff",
    x"00040000000001ffcd400000000000000000000000ff",
    x"00040000000000027fff0000000000000000000000ff",
    x"00040000000001b640000000000000000000000000ff",
    x"0004000000000107ffff0000000000000000000000ff",
    x"00040000000000006c1a0000000000000000000000ff",
    x"00040000000001e037c30000000000000000000000ff",
    x"00040000000001b6679f0000000000000000000000ff",
    x"00040000000001c904010000000000000000000000ff",
    x"000400000000003f7ff10000000000000000000000ff",
    x"000400000000000805e20000000000000000000000ff",
    x"00040000000000ff415c0000000000000000000000ff",
    x"000400000000000dd0ff0000000000000000000000ff",
    x"00040000000000e2f0100000000000000000000000ff",
    x"0004000000000194fbff0000000000000000000000ff",
    x"0004000000000099281a0000000000000000000000ff",
    x"00040000000001f1d6b50000000000000000000000ff",
    x"000400000000016c992e0000000000000000000000ff",
    x"0004000000000110b1fb0000000000000000000000ff",
    x"000400000000003c98c10000000000000000000000ff",
    x"0004000000000030855e0000000000000000000000ff",
    x"00040000000001a9b7620000000000000000000000ff",
    x"00040000000001d08da40000000000000000000000ff",
    x"0004000000000164743e0000000000000000000000ff",
    x"00040000000001fffc980000000000000000000000ff",
    x"0004000000000000341a0000000000000000000000ff",
    x"00040000000001fa38c30000000000000000000000ff",
    x"0004000000000075bf9f0000000000000000000000ff",
    x"000400000000016f04000000000000000000000000ff",
    x"00040000000000ff7ff10000000000000000000000ff",
    x"0004000000000008017c0000000000000000000000ff",
    x"00040000000000ffca610000000000000000000000ff",
    x"00040000000000014edf0000000000000000000000ff",
    x"00040000000001b938100000000000000000000000ff",
    x"000400000000002f7bff0000000000000000000000ff",
    x"0004000000000000101a0000000000000000000000ff",
    x"00040000000001fd8c000000000000000000000000ff",
    x"0004000000000040ffff0000000000000000000000ff",
    x"00040000000001b000000000000000000000000000ff",
    x"00040000000001fffff70000000000000000000000ff",
    x"000400000000000001820000000000000000000000ff",
    x"00040000000001ffcd400000000000000000000000ff",
    x"00040000000000027fff0000000000000000000000ff",
    x"00040000000001b640000000000000000000000000ff",
    x"0004000000000107ffff0000000000000000000000ff"
  );
end package;