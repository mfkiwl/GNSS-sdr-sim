library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package input is
  
  constant inputFrameSatCount : integer := 1;
  
  type inputTable is array(0 to 1810 - 1) of std_logic_vector(176-1 downto 0);
  constant inputSeq : inputTable := (
    x"ffff0000000000000011000001021fcd03fff5ecbbff",
    x"ffff000000000000000600000000001f1dfff5ecb1ff",
    x"ffff00000000000000000000000000288ffff5eca6ff",
    x"ffff00000000000000000000000000288efff5ec9bff",
    x"ffff00000000000000000000000000288ffff5ec91ff",
    x"ffff00000000000000090000000000288ffff5ec86ff",
    x"ffff000000000000000a00000000002890fff5ec7cff",
    x"ffff00000000000000110000000000288ffff5ec71ff",
    x"ffff000000000000000100000000002890fff5ec66ff",
    x"ffff00000000000000020000000000288ffff5ec5cff",
    x"ffff000000000000001600000000002890fff5ec51ff",
    x"ffff000000000000000600000000002890fff5ec47ff",
    x"ffff000000000000001c00000000002891fff5ec3cff",
    x"ffff000000000000001100000000002890fff5ec31ff",
    x"ffff000000000000000200000000002891fff5ec27ff",
    x"ffff000000000000000000000000002890fff5ec1cff",
    x"ffff000000000000001000000000002891fff5ec12ff",
    x"ffff000000000000000400000000002891fff5ec07ff",
    x"ffff000000000000000000000000002892fff5ebfdff",
    x"ffff000000000000000000000000002891fff5ebf2ff",
    x"ffff000000000000000000000000002892fff5ebe7ff",
    x"ffff000000000000000000000000002891fff5ebddff",
    x"ffff000000000000000000000000002892fff5ebd2ff",
    x"ffff000000000000000000000000002892fff5ebc8ff",
    x"ffff000000000000000000000000002893fff5ebbdff",
    x"ffff000000000000000000000000002892fff5ebb2ff",
    x"ffff000000000000000000000000002892fff5eba8ff",
    x"ffff000000000000000000000000002893fff5eb9dff",
    x"ffff000000000000000000000000002893fff5eb93ff",
    x"ffff000000000000000000000000002893fff5eb88ff",
    x"ffff000000000000000000000000002893fff5eb7dff",
    x"ffff000000000000000000000000002894fff5eb73ff",
    x"ffff000000000000000000000000002893fff5eb68ff",
    x"ffff000000000000000000000000002894fff5eb5eff",
    x"ffff000000000000000000000000002894fff5eb53ff",
    x"ffff000000000000000000000000002894fff5eb48ff",
    x"ffff000000000000000000000000002894fff5eb3eff",
    x"ffff000000000000000000000000002895fff5eb33ff",
    x"ffff000000000000000000000000002894fff5eb29ff",
    x"ffff000000000000000e00000000002895fff5eb1eff",
    x"ffff000000000000000100000000002895fff5eb14ff",
    x"ffff000000000000001b00000000002895fff5eb09ff",
    x"ffff000000000000000500000000002895fff5eafeff",
    x"ffff000000000000001900000000002896fff5eaf4ff",
    x"ffff000000000000001f00000000002895fff5eae9ff",
    x"ffff000000000000001f00000000002896fff5eadfff",
    x"ffff000000000000001f00000000002896fff5ead4ff",
    x"ffff000000000000001e00000000002896fff5eac9ff",
    x"ffff000000000000001f00000000002896fff5eabfff",
    x"ffff000000000000000700000000002897fff5eab4ff",
    x"ffff000000000000000000000000002896fff5eaaaff",
    x"ffff000000000000000000000000002897fff5ea9fff",
    x"ffff000000000000000300000000002897fff5ea94ff",
    x"ffff000000000000001d00000000002897fff5ea8aff",
    x"ffff000000000000000800000000002897fff5ea7fff",
    x"ffff000000000000001e00000000002897fff5ea75ff",
    x"ffff000000000000000a00000000002898fff5ea6aff",
    x"ffff000000000000000000000000002898fff5ea5fff",
    x"ffff000000000000001400000000002898fff5ea55ff",
    x"ffff000000000000000100000000002898fff5ea4aff",
    x"ffff000000000000001100000000002898fff5ea40ff",
    x"ffff000000000000000600000000002898fff5ea35ff",
    x"ffff000000000000000000000000002899fff5ea2bff",
    x"ffff000000000000000000000000002899fff5ea20ff",
    x"ffff000000000000000000000000002899fff5ea15ff",
    x"ffff000000000000000900000000002899fff5ea0bff",
    x"ffff000000000000000a00000000002899fff5ea00ff",
    x"ffff000000000000001100000000002899fff5e9f6ff",
    x"ffff00000000000000010000000000289afff5e9ebff",
    x"ffff00000000000000010000000000289afff5e9e0ff",
    x"ffff000000000000001100000000002899fff5e9d6ff",
    x"ffff00000000000000070000000000289bfff5e9cbff",
    x"ffff000000000000001a0000000000289afff5e9c1ff",
    x"ffff00000000000000060000000000289afff5e9b6ff",
    x"ffff00000000000000100000000000289bfff5e9abff",
    x"ffff00000000000000110000000000289afff5e9a1ff",
    x"ffff00000000000000190000000000289bfff5e996ff",
    x"ffff00000000000000020000000000289bfff5e98cff",
    x"ffff000000000000000c0000000000289cfff5e981ff",
    x"ffff00000000000000140000000000289bfff5e976ff",
    x"ffff000000000000001e0000000000289cfff5e96cff",
    x"ffff00000000000000180000000000289bfff5e961ff",
    x"ffff00000000000000160000000000289cfff5e957ff",
    x"ffff000000000000000d0000000000289cfff5e94cff",
    x"ffff00000000000000020000000000289dfff5e941ff",
    x"ffff00000000000000020000000000289cfff5e937ff",
    x"ffff00000000000000030000000000289dfff5e92cff",
    x"ffff00000000000000190000000000289cfff5e922ff",
    x"ffff00000000000000060000000000289dfff5e917ff",
    x"ffff000000000000001b0000000000289dfff5e90dff",
    x"ffff000000000000001f0000000000289dfff5e902ff",
    x"ffff000000000000000d0000000000289efff5e8f7ff",
    x"ffff00000000000000100000000000289dfff5e8edff",
    x"ffff000000000000001e0000000000289efff5e8e2ff",
    x"ffff00000000000000130000000000289efff5e8d8ff",
    x"ffff00000000000000050000000000289efff5e8cdff",
    x"ffff00000000000000000000000000289efff5e8c2ff",
    x"ffff00000000000000040000000000289ffff5e8b8ff",
    x"ffff000000000000001b0000000000289efff5e8adff",
    x"ffff00000000000000150000000000289ffff5e8a3ff",
    x"ffff00000000000000070000000000289ffff5e898ff",
    x"ffff00000000000000160000000000289ffff5e88dff",
    x"ffff000000000000000f0000000000289ffff5e883ff",
    x"ffff0000000000000001000000000028a0fff5e878ff",
    x"ffff00000000000000180000000000289ffff5e86eff",
    x"ffff0000000000000014000000000028a0fff5e863ff",
    x"ffff0000000000000007000000000028a0fff5e858ff",
    x"ffff0000000000000007000000000028a0fff5e84eff",
    x"ffff0000000000000010000000000028a0fff5e843ff",
    x"ffff0000000000000003000000000028a0fff5e839ff",
    x"ffff0000000000000012000000000028a1fff5e82eff",
    x"ffff000000000000001f000000000028a1fff5e823ff",
    x"ffff0000000000000001000000000028a1fff5e819ff",
    x"ffff0000000000000007000000000028a1fff5e80eff",
    x"ffff000000000000001c000000000028a1fff5e804ff",
    x"ffff0000000000000017000000000028a1fff5e7f9ff",
    x"ffff0000000000000004000000000028a2fff5e7eeff",
    x"ffff0000000000000000000000000028a2fff5e7e4ff",
    x"ffff000000000000000c000000000028a2fff5e7d9ff",
    x"ffff0000000000000000000000000028a5fff5e7cfff",
    x"ffff0000000000000011000000000028a2fff5e7c4ff",
    x"ffff0000000000000006000000000028a2fff5e7baff",
    x"ffff0000000000000000000000000028a3fff5e7afff",
    x"ffff0000000000000000000000000028a2fff5e7a4ff",
    x"ffff0000000000000000000000000028a3fff5e79aff",
    x"ffff0000000000000009000000000028a3fff5e78fff",
    x"ffff000000000000000a000000000028a4fff5e785ff",
    x"ffff0000000000000011000000000028a3fff5e77aff",
    x"ffff0000000000000001000000000028a4fff5e76fff",
    x"ffff0000000000000003000000000028a3fff5e765ff",
    x"ffff0000000000000017000000000028a4fff5e75aff",
    x"ffff0000000000000005000000000028a4fff5e750ff",
    x"ffff000000000000001f000000000028a5fff5e745ff",
    x"ffff000000000000001f000000000028a4fff5e73aff",
    x"ffff0000000000000002000000000028a4fff5e730ff",
    x"ffff0000000000000000000000000028a5fff5e725ff",
    x"ffff0000000000000012000000000028a5fff5e71bff",
    x"ffff0000000000000010000000000028a5fff5e710ff",
    x"ffff0000000000000018000000000028a5fff5e705ff",
    x"ffff000000000000001e000000000028a6fff5e6fbff",
    x"ffff0000000000000003000000000028a5fff5e6f0ff",
    x"ffff000000000000001f000000000028a6fff5e6e6ff",
    x"ffff000000000000000d000000000028a6fff5e6dbff",
    x"ffff0000000000000019000000000028a6fff5e6d0ff",
    x"ffff0000000000000000000000000028a6fff5e6c6ff",
    x"ffff0000000000000000000000000028a7fff5e6bbff",
    x"ffff0000000000000002000000000028a6fff5e6b1ff",
    x"ffff0000000000000016000000000028a7fff5e6a6ff",
    x"ffff0000000000000011000000000028a7fff5e69bff",
    x"ffff000000000000000a000000000028a7fff5e691ff",
    x"ffff000000000000001e000000000028a7fff5e686ff",
    x"ffff000000000000001c000000000028a7fff5e67cff",
    x"ffff000000000000001e000000000028a8fff5e671ff",
    x"ffff0000000000000004000000000028a8fff5e666ff",
    x"ffff0000000000000005000000000028a8fff5e65cff",
    x"ffff0000000000000013000000000028a8fff5e651ff",
    x"ffff000000000000001b000000000028a8fff5e647ff",
    x"ffff0000000000000005000000000028a8fff5e63cff",
    x"ffff000000000000000f000000000028a9fff5e631ff",
    x"ffff0000000000000006000000000028a9fff5e627ff",
    x"ffff000000000000000b000000000028a9fff5e61cff",
    x"ffff0000000000000009000000000028a9fff5e612ff",
    x"ffff0000000000000011000000000028a9fff5e607ff",
    x"ffff0000000000000003000000000028a9fff5e5fcff",
    x"ffff0000000000000018000000000028aafff5e5f2ff",
    x"ffff0000000000000002000000000028a9fff5e5e7ff",
    x"ffff0000000000000009000000000028aafff5e5ddff",
    x"ffff0000000000000018000000000028aafff5e5d2ff",
    x"ffff0000000000000000000000000028abfff5e5c7ff",
    x"ffff0000000000000010000000000028aafff5e5bdff",
    x"ffff0000000000000016000000000028abfff5e5b2ff",
    x"ffff0000000000000014000000000028aafff5e5a8ff",
    x"ffff0000000000000002000000000028abfff5e59dff",
    x"ffff0000000000000001000000000028abfff5e592ff",
    x"ffff000000000000001a000000000028abfff5e588ff",
    x"ffff0000000000000006000000000028acfff5e57dff",
    x"ffff0000000000000014000000000028abfff5e573ff",
    x"ffff000000000000001c000000000028acfff5e568ff",
    x"ffff0000000000000019000000000028acfff5e55dff",
    x"ffff0000000000000001000000000028acfff5e553ff",
    x"ffff0000000000000011000000000028acfff5e548ff",
    x"ffff0000000000000006000000000028adfff5e53eff",
    x"ffff0000000000000000000000000028acfff5e533ff",
    x"ffff0000000000000000000000000028adfff5e528ff",
    x"ffff0000000000000000000000000028adfff5e51eff",
    x"ffff0000000000000009000000000028adfff5e513ff",
    x"ffff000000000000000a000000000028adfff5e509ff",
    x"ffff0000000000000011000000000028aefff5e4feff",
    x"ffff0000000000000011000000000028adfff5e4f3ff",
    x"ffff0000000000000010000000000028aefff5e4e9ff",
    x"ffff0000000000000008000000000028aefff5e4deff",
    x"ffff0000000000000004000000000028aefff5e4d4ff",
    x"ffff000000000000001d000000000028aefff5e4c9ff",
    x"ffff0000000000000004000000000028aefff5e4beff",
    x"ffff0000000000000000000000000028affff5e4b4ff",
    x"ffff0000000000000000000000000028affff5e4a9ff",
    x"ffff0000000000000010000000000028affff5e49fff",
    x"ffff000000000000001e000000000028affff5e494ff",
    x"ffff000000000000001f000000000028affff5e489ff",
    x"ffff000000000000001f000000000028affff5e47fff",
    x"ffff000000000000001f000000000028b0fff5e474ff",
    x"ffff000000000000001f000000000028b0fff5e46aff",
    x"ffff000000000000001f000000000028b0fff5e45fff",
    x"ffff000000000000001f000000000028affff5e454ff",
    x"ffff000000000000001f000000000028b1fff5e44aff",
    x"ffff000000000000001f000000000028b0fff5e43fff",
    x"ffff000000000000001f000000000028b1fff5e435ff",
    x"ffff000000000000001f000000000028b0fff5e42aff",
    x"ffff000000000000001f000000000028b1fff5e41fff",
    x"ffff000000000000001f000000000028b1fff5e415ff",
    x"ffff000000000000001f000000000028b2fff5e40aff",
    x"ffff000000000000001f000000000028b1fff5e400ff",
    x"ffff000000000000001f000000000028b2fff5e3f5ff",
    x"ffff000000000000001f000000000028b1fff5e3eaff",
    x"ffff000000000000001f000000000028b2fff5e3e0ff",
    x"ffff000000000000001f000000000028b2fff5e3d5ff",
    x"ffff000000000000001f000000000028b2fff5e3cbff",
    x"ffff000000000000001f000000000028b3fff5e3c0ff",
    x"ffff000000000000001f000000000028b2fff5e3b5ff",
    x"ffff000000000000001f000000000028b3fff5e3abff",
    x"ffff000000000000001f000000000028b3fff5e3a0ff",
    x"ffff000000000000001f000000000028b3fff5e396ff",
    x"ffff000000000000001f000000000028b3fff5e38bff",
    x"ffff000000000000001f000000000028b4fff5e380ff",
    x"ffff000000000000001f000000000028b3fff5e376ff",
    x"ffff000000000000001f000000000028b4fff5e36bff",
    x"ffff000000000000001f000000000028b4fff5e361ff",
    x"ffff000000000000001f000000000028b4fff5e356ff",
    x"ffff000000000000001f000000000028b4fff5e34bff",
    x"ffff000000000000001f000000000028b5fff5e341ff",
    x"ffff000000000000001f000000000028b4fff5e336ff",
    x"ffff000000000000001f000000000028b5fff5e32cff",
    x"ffff000000000000001f000000000028b5fff5e321ff",
    x"ffff000000000000001f000000000028b5fff5e316ff",
    x"ffff000000000000001f000000000028b5fff5e30cff",
    x"ffff000000000000001f000000000028b5fff5e301ff",
    x"ffff000000000000001f000000000028b6fff5e2f7ff",
    x"ffff000000000000001f000000000028b6fff5e2ecff",
    x"ffff0000000000000017000000000028b6fff5e2e1ff",
    x"ffff0000000000000006000000000028b6fff5e2d7ff",
    x"ffff0000000000000011000000000028b6fff5e2ccff",
    x"ffff0000000000000006000000000028b6fff5e2c2ff",
    x"ffff0000000000000000000000000028b7fff5e2b7ff",
    x"ffff0000000000000000000000000028b7fff5e2acff",
    x"ffff0000000000000000000000000028b6fff5e2a2ff",
    x"ffff0000000000000009000000000028b8fff5e297ff",
    x"ffff000000000000000a000000000028b7fff5e28dff",
    x"ffff0000000000000011000000000028b7fff5e282ff",
    x"ffff0000000000000011000000000028b8fff5e277ff",
    x"ffff0000000000000012000000000028b7fff5e26dff",
    x"ffff000000000000000e000000000028b8fff5e262ff",
    x"ffff0000000000000006000000000028b8fff5e258ff",
    x"ffff0000000000000012000000000028b9fff5e24dff",
    x"ffff0000000000000010000000000028b8fff5e242ff",
    x"ffff0000000000000004000000000028b9fff5e238ff",
    x"ffff0000000000000005000000000028b8fff5e22dff",
    x"ffff000000000000000c000000000028b9fff5e223ff",
    x"ffff000000000000001e000000000028b9fff5e218ff",
    x"ffff000000000000001f000000000028b9fff5e20dff",
    x"ffff000000000000001b000000000028bafff5e203ff",
    x"ffff0000000000000009000000000028b9fff5e1f8ff",
    x"ffff0000000000000002000000000028bafff5e1eeff",
    x"ffff000000000000001e000000000028bafff5e1e3ff",
    x"ffff000000000000001d000000000028bafff5e1d8ff",
    x"ffff0000000000000010000000000028bafff5e1ceff",
    x"ffff0000000000000004000000000028bbfff5e1c3ff",
    x"ffff0000000000000006000000000028bafff5e1b8ff",
    x"ffff000000000000001f000000000028bbfff5e1aeff",
    x"ffff000000000000000f000000000028bbfff5e1a3ff",
    x"ffff000000000000001f000000000028bbfff5e199ff",
    x"ffff000000000000001a000000000028befff5e18eff",
    x"ffff000000000000001b000000000028bcfff5e183ff",
    x"ffff0000000000000003000000000028bbfff5e179ff",
    x"ffff000000000000001b000000000028bcfff5e16eff",
    x"ffff000000000000000f000000000028bcfff5e164ff",
    x"ffff0000000000000016000000000028bcfff5e159ff",
    x"ffff000000000000001f000000000028bcfff5e14eff",
    x"ffff000000000000000a000000000028bcfff5e144ff",
    x"ffff000000000000001a000000000028bdfff5e139ff",
    x"ffff0000000000000019000000000028bdfff5e12fff",
    x"ffff000000000000000f000000000028bdfff5e124ff",
    x"ffff000000000000001d000000000028bdfff5e119ff",
    x"ffff000000000000001b000000000028bdfff5e10fff",
    x"ffff0000000000000011000000000028bdfff5e104ff",
    x"ffff0000000000000003000000000028befff5e0faff",
    x"ffff000000000000001a000000000028befff5e0efff",
    x"ffff0000000000000014000000000028befff5e0e4ff",
    x"ffff000000000000000b000000000028befff5e0daff",
    x"ffff000000000000001e000000000028befff5e0cfff",
    x"ffff0000000000000009000000000028befff5e0c5ff",
    x"ffff0000000000000009000000000028bffff5e0baff",
    x"ffff000000000000001c000000000028bffff5e0afff",
    x"ffff000000000000001b000000000028befff5e0a5ff",
    x"ffff0000000000000018000000000028bffff5e09aff",
    x"ffff0000000000000008000000000028c0fff5e090ff",
    x"ffff0000000000000006000000000028bffff5e085ff",
    x"ffff0000000000000000000000000028c0fff5e07aff",
    x"ffff0000000000000000000000000028bffff5e070ff",
    x"ffff0000000000000018000000000028c0fff5e065ff",
    x"ffff0000000000000004000000000028c0fff5e05bff",
    x"ffff0000000000000011000000000028c1fff5e050ff",
    x"ffff0000000000000006000000000028c0fff5e045ff",
    x"ffff0000000000000000000000000028c0fff5e03bff",
    x"ffff0000000000000000000000000028c1fff5e030ff",
    x"ffff0000000000000000000000000028c1fff5e025ff",
    x"ffff0000000000000009000000000028c1fff5e01bff",
    x"ffff000000000000000a000000000028c2fff5e010ff",
    x"ffff0000000000000011000000000028c1fff5e006ff",
    x"ffff0000000000000011000000000028c1fff5dffbff",
    x"ffff0000000000000001000000000028c2fff5dff0ff",
    x"ffff000000000000000e000000000028c2fff5dfe6ff",
    x"ffff0000000000000002000000000028c2fff5dfdbff",
    x"ffff000000000000001c000000000028c2fff5dfd1ff",
    x"ffff0000000000000011000000000028c3fff5dfc6ff",
    x"ffff0000000000000002000000000028c2fff5dfbbff",
    x"ffff0000000000000000000000000028c3fff5dfb1ff",
    x"ffff0000000000000010000000000028c3fff5dfa6ff",
    x"ffff0000000000000004000000000028c3fff5df9cff",
    x"ffff0000000000000000000000000028c3fff5df91ff",
    x"ffff0000000000000000000000000028c4fff5df86ff",
    x"ffff0000000000000000000000000028c3fff5df7cff",
    x"ffff0000000000000000000000000028c4fff5df71ff",
    x"ffff0000000000000000000000000028c4fff5df67ff",
    x"ffff0000000000000000000000000028c4fff5df5cff",
    x"ffff0000000000000000000000000028c4fff5df51ff",
    x"ffff0000000000000000000000000028c5fff5df47ff",
    x"ffff0000000000000000000000000028c4fff5df3cff",
    x"ffff0000000000000000000000000028c5fff5df32ff",
    x"ffff0000000000000000000000000028c5fff5df27ff",
    x"ffff0000000000000000000000000028c5fff5df1cff",
    x"ffff0000000000000000000000000028c5fff5df12ff",
    x"ffff0000000000000000000000000028c5fff5df07ff",
    x"ffff0000000000000000000000000028c6fff5defcff",
    x"ffff0000000000000000000000000028c6fff5def2ff",
    x"ffff0000000000000000000000000028c6fff5dee7ff",
    x"ffff0000000000000000000000000028c6fff5deddff",
    x"ffff0000000000000000000000000028c6fff5ded2ff",
    x"ffff0000000000000000000000000028c6fff5dec7ff",
    x"ffff0000000000000000000000000028c7fff5debdff",
    x"ffff000000000000000e000000000028c7fff5deb2ff",
    x"ffff0000000000000001000000000028c7fff5dea8ff",
    x"ffff000000000000001b000000000028c7fff5de9dff",
    x"ffff0000000000000005000000000028c7fff5de92ff",
    x"ffff0000000000000019000000000028c7fff5de88ff",
    x"ffff000000000000001f000000000028c8fff5de7dff",
    x"ffff000000000000001f000000000028c8fff5de73ff",
    x"ffff000000000000001f000000000028c8fff5de68ff",
    x"ffff000000000000001e000000000028c8fff5de5dff",
    x"ffff000000000000001f000000000028c8fff5de53ff",
    x"ffff0000000000000007000000000028c8fff5de48ff",
    x"ffff0000000000000000000000000028c9fff5de3eff",
    x"ffff0000000000000000000000000028c9fff5de33ff",
    x"ffff0000000000000003000000000028c8fff5de28ff",
    x"ffff000000000000001d000000000028cafff5de1eff",
    x"ffff0000000000000008000000000028c9fff5de13ff",
    x"ffff000000000000001e000000000028c9fff5de08ff",
    x"ffff000000000000000a000000000028cafff5ddfeff",
    x"ffff0000000000000000000000000028c9fff5ddf3ff",
    x"ffff0000000000000014000000000028cafff5dde9ff",
    x"ffff0000000000000001000000000028cafff5dddeff",
    x"ffff0000000000000011000000000028cbfff5ddd3ff",
    x"ffff0000000000000006000000000028cafff5ddc9ff",
    x"ffff0000000000000000000000000028cbfff5ddbeff",
    x"ffff0000000000000000000000000028cafff5ddb4ff",
    x"ffff0000000000000000000000000028cbfff5dda9ff",
    x"ffff0000000000000009000000000028cbfff5dd9eff",
    x"ffff000000000000000a000000000028ccfff5dd94ff",
    x"ffff0000000000000011000000000028cbfff5dd89ff",
    x"ffff0000000000000011000000000028ccfff5dd7fff",
    x"ffff0000000000000003000000000028cbfff5dd74ff",
    x"ffff0000000000000015000000000028ccfff5dd69ff",
    x"ffff0000000000000000000000000028ccfff5dd5fff",
    x"ffff000000000000001a000000000028cdfff5dd54ff",
    x"ffff0000000000000006000000000028ccfff5dd49ff",
    x"ffff0000000000000010000000000028cdfff5dd3fff",
    x"ffff0000000000000011000000000028ccfff5dd34ff",
    x"ffff0000000000000019000000000028cdfff5dd2aff",
    x"ffff0000000000000002000000000028cdfff5dd1fff",
    x"ffff000000000000000c000000000028cefff5dd14ff",
    x"ffff0000000000000014000000000028cdfff5dd0aff",
    x"ffff000000000000001e000000000028cdfff5dcffff",
    x"ffff0000000000000018000000000028cefff5dcf5ff",
    x"ffff0000000000000016000000000028cefff5dceaff",
    x"ffff000000000000000d000000000028cefff5dcdfff",
    x"ffff0000000000000002000000000028cefff5dcd5ff",
    x"ffff0000000000000002000000000028cffff5dccaff",
    x"ffff0000000000000003000000000028cefff5dcc0ff",
    x"ffff0000000000000019000000000028cffff5dcb5ff",
    x"ffff0000000000000006000000000028cffff5dcaaff",
    x"ffff000000000000001b000000000028cffff5dca0ff",
    x"ffff000000000000001f000000000028cffff5dc95ff",
    x"ffff000000000000000d000000000028d0fff5dc8aff",
    x"ffff0000000000000010000000000028cffff5dc80ff",
    x"ffff000000000000001e000000000028d0fff5dc75ff",
    x"ffff0000000000000013000000000028d0fff5dc6bff",
    x"ffff0000000000000005000000000028d0fff5dc60ff",
    x"ffff0000000000000000000000000028d0fff5dc55ff",
    x"ffff0000000000000004000000000028d1fff5dc4bff",
    x"ffff000000000000001b000000000028d0fff5dc40ff",
    x"ffff0000000000000015000000000028d1fff5dc36ff",
    x"ffff0000000000000007000000000028d1fff5dc2bff",
    x"ffff0000000000000016000000000028d1fff5dc20ff",
    x"ffff000000000000000f000000000028d1fff5dc16ff",
    x"ffff0000000000000001000000000028d2fff5dc0bff",
    x"ffff0000000000000018000000000028d1fff5dc01ff",
    x"ffff0000000000000014000000000028d2fff5dbf6ff",
    x"ffff0000000000000007000000000028d2fff5dbebff",
    x"ffff0000000000000007000000000028d2fff5dbe1ff",
    x"ffff0000000000000010000000000028d2fff5dbd6ff",
    x"ffff0000000000000003000000000028d3fff5dbcbff",
    x"ffff0000000000000012000000000028d2fff5dbc1ff",
    x"ffff000000000000001f000000000028d3fff5dbb6ff",
    x"ffff0000000000000001000000000028d3fff5dbacff",
    x"ffff0000000000000007000000000028d3fff5dba1ff",
    x"ffff000000000000001c000000000028d3fff5db96ff",
    x"ffff0000000000000017000000000028d4fff5db8cff",
    x"ffff0000000000000004000000000028d3fff5db81ff",
    x"ffff0000000000000000000000000028d4fff5db77ff",
    x"ffff000000000000000c000000000028d4fff5db6cff",
    x"ffff0000000000000000000000000028d4fff5db61ff",
    x"ffff0000000000000011000000000028d4fff5db57ff",
    x"ffff0000000000000006000000000028d8fff5db4cff",
    x"ffff0000000000000000000000000028d4fff5db41ff",
    x"ffff0000000000000000000000000028d5fff5db37ff",
    x"ffff0000000000000000000000000028d5fff5db2cff",
    x"ffff0000000000000009000000000028d5fff5db22ff",
    x"ffff000000000000000a000000000028d5fff5db17ff",
    x"ffff0000000000000011000000000028d6fff5db0cff",
    x"ffff0000000000000009000000000028d5fff5db02ff",
    x"ffff0000000000000000000000000028d6fff5daf7ff",
    x"ffff000000000000000b000000000028d6fff5daedff",
    x"ffff0000000000000005000000000028d6fff5dae2ff",
    x"ffff000000000000001f000000000028d6fff5dad7ff",
    x"ffff000000000000001f000000000028d7fff5dacdff",
    x"ffff0000000000000002000000000028d6fff5dac2ff",
    x"ffff0000000000000000000000000028d7fff5dab7ff",
    x"ffff0000000000000012000000000028d7fff5daadff",
    x"ffff0000000000000010000000000028d7fff5daa2ff",
    x"ffff0000000000000018000000000028d7fff5da98ff",
    x"ffff000000000000001e000000000028d8fff5da8dff",
    x"ffff0000000000000003000000000028d7fff5da82ff",
    x"ffff000000000000001f000000000028d8fff5da78ff",
    x"ffff000000000000000d000000000028d8fff5da6dff",
    x"ffff0000000000000019000000000028d8fff5da63ff",
    x"ffff0000000000000000000000000028d8fff5da58ff",
    x"ffff0000000000000000000000000028d9fff5da4dff",
    x"ffff0000000000000002000000000028d9fff5da43ff",
    x"ffff0000000000000016000000000028d8fff5da38ff",
    x"ffff0000000000000011000000000028d9fff5da2dff",
    x"ffff000000000000000a000000000028d9fff5da23ff",
    x"ffff000000000000001e000000000028dafff5da18ff",
    x"ffff000000000000001c000000000028d9fff5da0eff",
    x"ffff000000000000001e000000000028dafff5da03ff",
    x"ffff0000000000000004000000000028d9fff5d9f8ff",
    x"ffff0000000000000005000000000028dafff5d9eeff",
    x"ffff0000000000000013000000000028dafff5d9e3ff",
    x"ffff000000000000001b000000000028dbfff5d9d9ff",
    x"ffff0000000000000005000000000028dafff5d9ceff",
    x"ffff000000000000000f000000000028dbfff5d9c3ff",
    x"ffff0000000000000006000000000028dafff5d9b9ff",
    x"ffff000000000000000b000000000028dbfff5d9aeff",
    x"ffff0000000000000009000000000028dbfff5d9a4ff",
    x"ffff0000000000000011000000000028dcfff5d999ff",
    x"ffff0000000000000003000000000028dbfff5d98eff",
    x"ffff0000000000000018000000000028dcfff5d984ff",
    x"ffff0000000000000002000000000028dbfff5d979ff",
    x"ffff0000000000000009000000000028dcfff5d96eff",
    x"ffff0000000000000018000000000028dcfff5d964ff",
    x"ffff0000000000000000000000000028ddfff5d959ff",
    x"ffff0000000000000010000000000028dcfff5d94fff",
    x"ffff0000000000000016000000000028ddfff5d944ff",
    x"ffff0000000000000014000000000028ddfff5d939ff",
    x"ffff0000000000000002000000000028dcfff5d92fff",
    x"ffff0000000000000001000000000028defff5d924ff",
    x"ffff000000000000001a000000000028ddfff5d919ff",
    x"ffff0000000000000006000000000028ddfff5d90fff",
    x"ffff0000000000000014000000000028defff5d904ff",
    x"ffff000000000000001c000000000028defff5d8faff",
    x"ffff0000000000000019000000000028ddfff5d8efff",
    x"ffff0000000000000001000000000028dffff5d8e4ff",
    x"ffff0000000000000011000000000028defff5d8daff",
    x"ffff0000000000000006000000000028defff5d8cfff",
    x"ffff0000000000000000000000000028dffff5d8c5ff",
    x"ffff0000000000000000000000000028dffff5d8baff",
    x"ffff0000000000000000000000000028dffff5d8afff",
    x"ffff0000000000000009000000000028dffff5d8a5ff",
    x"ffff000000000000000a000000000028dffff5d89aff",
    x"ffff0000000000000011000000000028dffff5d88fff",
    x"ffff0000000000000009000000000028e0fff5d885ff",
    x"ffff0000000000000012000000000028e0fff5d87aff",
    x"ffff0000000000000000000000000028e0fff5d870ff",
    x"ffff0000000000000001000000000028e0fff5d865ff",
    x"ffff000000000000001d000000000028e0fff5d85aff",
    x"ffff0000000000000004000000000028e0fff5d850ff",
    x"ffff0000000000000000000000000028e1fff5d845ff",
    x"ffff0000000000000000000000000028e1fff5d83bff",
    x"ffff0000000000000010000000000028e1fff5d830ff",
    x"ffff000000000000001e000000000028e1fff5d825ff",
    x"ffff000000000000001f000000000028e1fff5d81bff",
    x"ffff000000000000001f000000000028e2fff5d810ff",
    x"ffff000000000000001f000000000028e1fff5d805ff",
    x"ffff000000000000001f000000000028e2fff5d7fbff",
    x"ffff000000000000001f000000000028e2fff5d7f0ff",
    x"ffff000000000000001f000000000028e2fff5d7e6ff",
    x"ffff000000000000001f000000000028e2fff5d7dbff",
    x"ffff000000000000001f000000000028e3fff5d7d0ff",
    x"ffff000000000000001f000000000028e2fff5d7c6ff",
    x"ffff000000000000001f000000000028e3fff5d7bbff",
    x"ffff000000000000001f000000000028e3fff5d7b0ff",
    x"ffff000000000000001f000000000028e3fff5d7a6ff",
    x"ffff000000000000001f000000000028e4fff5d79bff",
    x"ffff000000000000001f000000000028e3fff5d791ff",
    x"ffff000000000000001f000000000028e4fff5d786ff",
    x"ffff000000000000001f000000000028e3fff5d77bff",
    x"ffff000000000000001f000000000028e4fff5d771ff",
    x"ffff000000000000001f000000000028e4fff5d766ff",
    x"ffff000000000000001f000000000028e5fff5d75cff",
    x"ffff000000000000001f000000000028e4fff5d751ff",
    x"ffff000000000000001f000000000028e5fff5d746ff",
    x"ffff000000000000001f000000000028e4fff5d73cff",
    x"ffff000000000000001f000000000028e5fff5d731ff",
    x"ffff000000000000001f000000000028e6fff5d726ff",
    x"ffff000000000000001f000000000028e5fff5d71cff",
    x"ffff000000000000001f000000000028e5fff5d711ff",
    x"ffff000000000000001f000000000028e6fff5d707ff",
    x"ffff000000000000001f000000000028e6fff5d6fcff",
    x"ffff000000000000001f000000000028e6fff5d6f1ff",
    x"ffff000000000000001f000000000028e6fff5d6e7ff",
    x"ffff000000000000001f000000000028e6fff5d6dcff",
    x"ffff000000000000001f000000000028e6fff5d6d1ff",
    x"ffff000000000000001f000000000028e7fff5d6c7ff",
    x"ffff000000000000001f000000000028e7fff5d6bcff",
    x"ffff000000000000001f000000000028e7fff5d6b2ff",
    x"ffff000000000000001f000000000028e7fff5d6a7ff",
    x"ffff000000000000001f000000000028e7fff5d69cff",
    x"ffff000000000000001f000000000028e8fff5d692ff",
    x"ffff000000000000001f000000000028e7fff5d687ff",
    x"ffff000000000000001f000000000028e8fff5d67dff",
    x"ffff0000000000000017000000000028e8fff5d672ff",
    x"ffff0000000000000006000000000028e8fff5d667ff",
    x"ffff0000000000000011000000000028e8fff5d65dff",
    x"ffff0000000000000006000000000028e9fff5d652ff",
    x"ffff0000000000000000000000000028e8fff5d647ff",
    x"ffff0000000000000000000000000028e9fff5d63dff",
    x"ffff0000000000000000000000000028e9fff5d632ff",
    x"ffff0000000000000009000000000028e9fff5d628ff",
    x"ffff000000000000000a000000000028eafff5d61dff",
    x"ffff0000000000000011000000000028e9fff5d612ff",
    x"ffff0000000000000009000000000028eafff5d608ff",
    x"ffff0000000000000011000000000028e9fff5d5fdff",
    x"ffff000000000000001a000000000028eafff5d5f2ff",
    x"ffff0000000000000000000000000028ebfff5d5e8ff",
    x"ffff000000000000000a000000000028eafff5d5ddff",
    x"ffff0000000000000002000000000028eafff5d5d3ff",
    x"ffff000000000000001e000000000028ebfff5d5c8ff",
    x"ffff000000000000001d000000000028ebfff5d5bdff",
    x"ffff0000000000000000000000000028ebfff5d5b3ff",
    x"ffff000000000000001f000000000028ebfff5d5a8ff",
    x"ffff000000000000001f000000000028ebfff5d59dff",
    x"ffff000000000000000b000000000028ecfff5d593ff",
    x"ffff000000000000001f000000000028ebfff5d588ff",
    x"ffff0000000000000012000000000028ecfff5d57eff",
    x"ffff000000000000001e000000000028ecfff5d573ff",
    x"ffff0000000000000008000000000028ecfff5d568ff",
    x"ffff000000000000000f000000000028ecfff5d55eff",
    x"ffff000000000000000f000000000028edfff5d553ff",
    x"ffff000000000000001a000000000028ecfff5d548ff",
    x"ffff0000000000000001000000000028edfff5d53eff",
    x"ffff0000000000000010000000000028edfff5d533ff",
    x"ffff0000000000000000000000000028edfff5d529ff",
    x"ffff0000000000000005000000000028eefff5d51eff",
    x"ffff0000000000000004000000000028edfff5d513ff",
    x"ffff000000000000000c000000000028eefff5d509ff",
    x"ffff0000000000000019000000000028f0fff5d4feff",
    x"ffff0000000000000010000000000028eefff5d4f3ff",
    x"ffff0000000000000004000000000028effff5d4e9ff",
    x"ffff0000000000000009000000000028eefff5d4deff",
    x"ffff000000000000000c000000000028eefff5d4d4ff",
    x"ffff000000000000000f000000000028effff5d4c9ff",
    x"ffff000000000000000b000000000028effff5d4beff",
    x"ffff0000000000000000000000000028effff5d4b4ff",
    x"ffff000000000000001c000000000028effff5d4a9ff",
    x"ffff0000000000000001000000000028effff5d49eff",
    x"ffff0000000000000005000000000028f0fff5d494ff",
    x"ffff000000000000001c000000000028effff5d489ff",
    x"ffff0000000000000012000000000028f0fff5d47fff",
    x"ffff0000000000000005000000000028f0fff5d474ff",
    x"ffff0000000000000012000000000028f0fff5d469ff",
    x"ffff0000000000000001000000000028f0fff5d45fff",
    x"ffff0000000000000017000000000028f1fff5d454ff",
    x"ffff0000000000000008000000000028f1fff5d449ff",
    x"ffff0000000000000006000000000028f0fff5d43fff",
    x"ffff000000000000001c000000000028f1fff5d434ff",
    x"ffff0000000000000000000000000028f1fff5d42aff",
    x"ffff0000000000000003000000000028f2fff5d41fff",
    x"ffff0000000000000018000000000028f1fff5d414ff",
    x"ffff000000000000001f000000000028f2fff5d40aff",
    x"ffff000000000000000b000000000028f2fff5d3ffff",
    x"ffff000000000000000b000000000028f2fff5d3f5ff",
    x"ffff0000000000000001000000000028f2fff5d3eaff",
    x"ffff0000000000000011000000000028f2fff5d3dfff",
    x"ffff0000000000000006000000000028f3fff5d3d5ff",
    x"ffff0000000000000000000000000028f2fff5d3caff",
    x"ffff0000000000000000000000000028f3fff5d3bfff",
    x"ffff0000000000000000000000000028f3fff5d3b5ff",
    x"ffff0000000000000009000000000028f3fff5d3aaff",
    x"ffff000000000000000a000000000028f3fff5d3a0ff",
    x"ffff0000000000000011000000000028f4fff5d395ff",
    x"ffff0000000000000009000000000028f4fff5d38aff",
    x"ffff0000000000000003000000000028f3fff5d380ff",
    x"ffff0000000000000006000000000028f4fff5d375ff",
    x"ffff0000000000000007000000000028f5fff5d36aff",
    x"ffff000000000000001c000000000028f4fff5d360ff",
    x"ffff0000000000000011000000000028f4fff5d355ff",
    x"ffff0000000000000002000000000028f5fff5d34bff",
    x"ffff0000000000000000000000000028f5fff5d340ff",
    x"ffff0000000000000010000000000028f5fff5d335ff",
    x"ffff0000000000000004000000000028f5fff5d32bff",
    x"ffff0000000000000000000000000028f5fff5d320ff",
    x"ffff0000000000000000000000000028f6fff5d315ff",
    x"ffff0000000000000000000000000028f5fff5d30bff",
    x"ffff0000000000000000000000000028f6fff5d300ff",
    x"ffff0000000000000000000000000028f6fff5d2f6ff",
    x"ffff0000000000000000000000000028f6fff5d2ebff",
    x"ffff0000000000000000000000000028f7fff5d2e0ff",
    x"ffff0000000000000000000000000028f6fff5d2d6ff",
    x"ffff0000000000000000000000000028f7fff5d2cbff",
    x"ffff0000000000000000000000000028f7fff5d2c0ff",
    x"ffff0000000000000000000000000028f6fff5d2b6ff",
    x"ffff0000000000000000000000000028f8fff5d2abff",
    x"ffff0000000000000000000000000028f7fff5d2a0ff",
    x"ffff0000000000000000000000000028f8fff5d296ff",
    x"ffff0000000000000000000000000028f7fff5d28bff",
    x"ffff0000000000000000000000000028f8fff5d281ff",
    x"ffff0000000000000000000000000028f8fff5d276ff",
    x"ffff0000000000000000000000000028f8fff5d26bff",
    x"ffff0000000000000000000000000028f8fff5d261ff",
    x"ffff0000000000000000000000000028f9fff5d256ff",
    x"ffff0000000000000000000000000028f9fff5d24cff",
    x"ffff000000000000000e000000000028f8fff5d241ff",
    x"ffff0000000000000001000000000028f9fff5d236ff",
    x"ffff000000000000001b000000000028fafff5d22cff",
    x"ffff0000000000000005000000000028f9fff5d221ff",
    x"ffff0000000000000019000000000028f9fff5d216ff",
    x"ffff000000000000001f000000000028fafff5d20cff",
    x"ffff000000000000001f000000000028fafff5d201ff",
    x"ffff000000000000001f000000000028fafff5d1f6ff",
    x"ffff000000000000001e000000000028fafff5d1ecff",
    x"ffff000000000000001f000000000028fafff5d1e1ff",
    x"ffff0000000000000007000000000028fbfff5d1d7ff",
    x"ffff0000000000000000000000000028fafff5d1ccff",
    x"ffff0000000000000000000000000028fbfff5d1c1ff",
    x"ffff0000000000000003000000000028fbfff5d1b7ff",
    x"ffff000000000000001d000000000028fcfff5d1acff",
    x"ffff0000000000000008000000000028fbfff5d1a1ff",
    x"ffff000000000000001e000000000028fbfff5d197ff",
    x"ffff000000000000000a000000000028fcfff5d18cff",
    x"ffff0000000000000000000000000028fcfff5d182ff",
    x"ffff0000000000000014000000000028fcfff5d177ff",
    x"ffff0000000000000001000000000028fcfff5d16cff",
    x"ffff0000000000000011000000000028fcfff5d162ff",
    x"ffff0000000000000006000000000028fdfff5d157ff",
    x"ffff0000000000000000000000000028fcfff5d14cff",
    x"ffff0000000000000000000000000028fdfff5d142ff",
    x"ffff0000000000000000000000000028fdfff5d137ff",
    x"ffff0000000000000009000000000028fdfff5d12dff",
    x"ffff000000000000000a000000000028fefff5d122ff",
    x"ffff0000000000000011000000000028fdfff5d117ff",
    x"ffff0000000000000019000000000028fefff5d10dff",
    x"ffff0000000000000000000000000028fefff5d102ff",
    x"ffff0000000000000009000000000028fefff5d0f7ff",
    x"ffff0000000000000000000000000028fefff5d0edff",
    x"ffff000000000000001a000000000028fefff5d0e2ff",
    x"ffff0000000000000006000000000028fffff5d0d8ff",
    x"ffff0000000000000010000000000028fefff5d0cdff",
    x"ffff0000000000000011000000000028fffff5d0c2ff",
    x"ffff0000000000000019000000000028fffff5d0b8ff",
    x"ffff0000000000000002000000000028fffff5d0adff",
    x"ffff000000000000000c00000000002900fff5d0a2ff",
    x"ffff0000000000000014000000000028fffff5d098ff",
    x"ffff000000000000001e00000000002900fff5d08dff",
    x"ffff000000000000001800000000002900fff5d083ff",
    x"ffff000000000000001600000000002900fff5d078ff",
    x"ffff000000000000000d00000000002900fff5d06dff",
    x"ffff000000000000000200000000002900fff5d063ff",
    x"ffff000000000000000200000000002901fff5d058ff",
    x"ffff000000000000000300000000002901fff5d04dff",
    x"ffff000000000000001900000000002900fff5d043ff",
    x"ffff000000000000000600000000002901fff5d038ff",
    x"ffff000000000000001b00000000002902fff5d02dff",
    x"ffff000000000000001f00000000002901fff5d023ff",
    x"ffff000000000000000d00000000002901fff5d018ff",
    x"ffff000000000000001000000000002902fff5d00eff",
    x"ffff000000000000001e00000000002902fff5d003ff",
    x"ffff000000000000001300000000002902fff5cff8ff",
    x"ffff000000000000000500000000002902fff5cfeeff",
    x"ffff000000000000000000000000002902fff5cfe3ff",
    x"ffff000000000000000400000000002903fff5cfd8ff",
    x"ffff000000000000001b00000000002903fff5cfceff",
    x"ffff000000000000001500000000002903fff5cfc3ff",
    x"ffff000000000000000700000000002903fff5cfb9ff",
    x"ffff000000000000001600000000002903fff5cfaeff",
    x"ffff000000000000000f00000000002903fff5cfa3ff",
    x"ffff000000000000000100000000002904fff5cf99ff",
    x"ffff000000000000001800000000002903fff5cf8eff",
    x"ffff000000000000001400000000002904fff5cf83ff",
    x"ffff000000000000000700000000002904fff5cf79ff",
    x"ffff000000000000000700000000002904fff5cf6eff",
    x"ffff000000000000001000000000002905fff5cf63ff",
    x"ffff000000000000000300000000002904fff5cf59ff",
    x"ffff000000000000001200000000002905fff5cf4eff",
    x"ffff000000000000001f00000000002905fff5cf44ff",
    x"ffff000000000000000100000000002905fff5cf39ff",
    x"ffff000000000000000700000000002905fff5cf2eff",
    x"ffff000000000000001c00000000002905fff5cf24ff",
    x"ffff000000000000001700000000002906fff5cf19ff",
    x"ffff000000000000000400000000002906fff5cf0eff",
    x"ffff000000000000000000000000002905fff5cf04ff",
    x"ffff000000000000000c00000000002906fff5cef9ff",
    x"ffff000000000000000000000000002907fff5ceefff",
    x"ffff000000000000001100000000002906fff5cee4ff",
    x"ffff000000000000000600000000002907fff5ced9ff",
    x"ffff000000000000000000000000002906fff5cecfff",
    x"ffff000000000000000000000000002907fff5cec4ff",
    x"ffff000000000000000000000000002907fff5ceb9ff",
    x"ffff00000000000000090000000000290afff5ceafff",
    x"ffff000000000000000a00000000002908fff5cea4ff",
    x"ffff000000000000001100000000002907fff5ce99ff",
    x"ffff000000000000001900000000002908fff5ce8fff",
    x"ffff000000000000000200000000002908fff5ce84ff",
    x"ffff000000000000000f00000000002908fff5ce7aff",
    x"ffff000000000000000200000000002908fff5ce6fff",
    x"ffff000000000000001f00000000002908fff5ce64ff",
    x"ffff000000000000001f00000000002909fff5ce5aff",
    x"ffff000000000000000200000000002909fff5ce4fff",
    x"ffff000000000000000000000000002908fff5ce44ff",
    x"ffff00000000000000120000000000290afff5ce3aff",
    x"ffff000000000000001000000000002909fff5ce2fff",
    x"ffff000000000000001800000000002909fff5ce25ff",
    x"ffff000000000000001e0000000000290afff5ce1aff",
    x"ffff000000000000000300000000002909fff5ce0fff",
    x"ffff000000000000001f0000000000290afff5ce05ff",
    x"ffff000000000000000d0000000000290afff5cdfaff",
    x"ffff00000000000000190000000000290afff5cdefff",
    x"ffff00000000000000000000000000290bfff5cde5ff",
    x"ffff00000000000000000000000000290afff5cddaff",
    x"ffff00000000000000020000000000290bfff5cdcfff",
    x"ffff00000000000000160000000000290bfff5cdc5ff",
    x"ffff00000000000000110000000000290bfff5cdbaff",
    x"ffff000000000000000a0000000000290bfff5cdb0ff",
    x"ffff000000000000001e0000000000290cfff5cda5ff",
    x"ffff000000000000001c0000000000290bfff5cd9aff",
    x"ffff000000000000001e0000000000290cfff5cd90ff",
    x"ffff00000000000000040000000000290cfff5cd85ff",
    x"ffff00000000000000050000000000290cfff5cd7aff",
    x"ffff00000000000000130000000000290cfff5cd70ff",
    x"ffff000000000000001b0000000000290cfff5cd65ff",
    x"ffff00000000000000050000000000290dfff5cd5aff",
    x"ffff000000000000000f0000000000290dfff5cd50ff",
    x"ffff00000000000000060000000000290cfff5cd45ff",
    x"ffff000000000000000b0000000000290efff5cd3bff",
    x"ffff00000000000000090000000000290dfff5cd30ff",
    x"ffff00000000000000110000000000290dfff5cd25ff",
    x"ffff00000000000000030000000000290efff5cd1bff",
    x"ffff00000000000000180000000000290dfff5cd10ff",
    x"ffff00000000000000020000000000290efff5cd05ff",
    x"ffff00000000000000090000000000290efff5ccfbff",
    x"ffff00000000000000180000000000290ffff5ccf0ff",
    x"ffff00000000000000000000000000290efff5cce6ff",
    x"ffff00000000000000100000000000290efff5ccdbff",
    x"ffff00000000000000160000000000290ffff5ccd0ff",
    x"ffff00000000000000140000000000290ffff5ccc6ff",
    x"ffff00000000000000020000000000290ffff5ccbbff",
    x"ffff00000000000000010000000000290ffff5ccb0ff",
    x"ffff000000000000001a00000000002910fff5cca6ff",
    x"ffff00000000000000060000000000290ffff5cc9bff",
    x"ffff000000000000001400000000002910fff5cc90ff",
    x"ffff000000000000001c00000000002910fff5cc86ff",
    x"ffff000000000000001900000000002910fff5cc7bff",
    x"ffff000000000000000100000000002910fff5cc71ff",
    x"ffff000000000000001100000000002911fff5cc66ff",
    x"ffff000000000000000600000000002910fff5cc5bff",
    x"ffff000000000000000000000000002911fff5cc51ff",
    x"ffff000000000000000000000000002911fff5cc46ff",
    x"ffff000000000000000000000000002911fff5cc3bff",
    x"ffff000000000000000900000000002911fff5cc31ff",
    x"ffff000000000000000a00000000002911fff5cc26ff",
    x"ffff000000000000001100000000002912fff5cc1bff",
    x"ffff000000000000001900000000002912fff5cc11ff",
    x"ffff000000000000001100000000002912fff5cc06ff",
    x"ffff000000000000001800000000002912fff5cbfcff",
    x"ffff000000000000000500000000002912fff5cbf1ff",
    x"ffff000000000000001d00000000002912fff5cbe6ff",
    x"ffff000000000000000400000000002913fff5cbdcff",
    x"ffff000000000000000000000000002913fff5cbd1ff",
    x"ffff000000000000000000000000002913fff5cbc6ff",
    x"ffff000000000000001000000000002913fff5cbbcff",
    x"ffff000000000000001e00000000002913fff5cbb1ff",
    x"ffff000000000000001f00000000002913fff5cba6ff",
    x"ffff000000000000001f00000000002914fff5cb9cff",
    x"ffff000000000000001f00000000002914fff5cb91ff",
    x"ffff000000000000001f00000000002913fff5cb87ff",
    x"ffff000000000000001f00000000002915fff5cb7cff",
    x"ffff000000000000001f00000000002914fff5cb71ff",
    x"ffff000000000000001f00000000002914fff5cb67ff",
    x"ffff000000000000001f00000000002915fff5cb5cff",
    x"ffff000000000000001f00000000002914fff5cb51ff",
    x"ffff000000000000001f00000000002915fff5cb47ff",
    x"ffff000000000000001f00000000002915fff5cb3cff",
    x"ffff000000000000001f00000000002916fff5cb31ff",
    x"ffff000000000000001f00000000002915fff5cb27ff",
    x"ffff000000000000001f00000000002916fff5cb1cff",
    x"ffff000000000000001f00000000002915fff5cb12ff",
    x"ffff000000000000001f00000000002916fff5cb07ff",
    x"ffff000000000000001f00000000002916fff5cafcff",
    x"ffff000000000000001f00000000002917fff5caf2ff",
    x"ffff000000000000001f00000000002916fff5cae7ff",
    x"ffff000000000000001f00000000002917fff5cadcff",
    x"ffff000000000000001f00000000002916fff5cad2ff",
    x"ffff000000000000001f00000000002917fff5cac7ff",
    x"ffff000000000000001f00000000002917fff5cabcff",
    x"ffff000000000000001f00000000002918fff5cab2ff",
    x"ffff000000000000001f00000000002917fff5caa7ff",
    x"ffff000000000000001f00000000002918fff5ca9dff",
    x"ffff000000000000001f00000000002917fff5ca92ff",
    x"ffff000000000000001f00000000002918fff5ca87ff",
    x"ffff000000000000001f00000000002918fff5ca7dff",
    x"ffff000000000000001f00000000002919fff5ca72ff",
    x"ffff000000000000001f00000000002918fff5ca67ff",
    x"ffff000000000000001f00000000002919fff5ca5dff",
    x"ffff000000000000001f00000000002918fff5ca52ff",
    x"ffff000000000000001f00000000002919fff5ca47ff",
    x"ffff000000000000001f00000000002919fff5ca3dff",
    x"ffff000000000000001f0000000000291afff5ca32ff",
    x"ffff000000000000001f00000000002919fff5ca27ff",
    x"ffff000000000000001f0000000000291afff5ca1dff",
    x"ffff000000000000001f00000000002919fff5ca12ff",
    x"ffff000000000000001f0000000000291afff5ca08ff",
    x"ffff00000000000000170000000000291bfff5c9fdff",
    x"ffff00000000000000060000000000291afff5c9f2ff",
    x"ffff00000000000000110000000000291afff5c9e8ff",
    x"ffff00000000000000060000000000291bfff5c9ddff",
    x"ffff00000000000000000000000000291afff5c9d2ff",
    x"ffff00000000000000000000000000291bfff5c9c8ff",
    x"ffff00000000000000000000000000291cfff5c9bdff",
    x"ffff00000000000000090000000000291bfff5c9b3ff",
    x"ffff000000000000000a0000000000291bfff5c9a8ff",
    x"ffff00000000000000110000000000291cfff5c99dff",
    x"ffff00000000000000190000000000291cfff5c993ff",
    x"ffff00000000000000130000000000291bfff5c988ff",
    x"ffff000000000000001e0000000000291dfff5c97dff",
    x"ffff00000000000000070000000000291cfff5c973ff",
    x"ffff00000000000000020000000000291cfff5c968ff",
    x"ffff00000000000000060000000000291dfff5c95dff",
    x"ffff00000000000000050000000000291dfff5c953ff",
    x"ffff00000000000000030000000000291dfff5c948ff",
    x"ffff000000000000000a0000000000291dfff5c93dff",
    x"ffff000000000000001f0000000000291dfff5c933ff",
    x"ffff000000000000001f0000000000291dfff5c928ff",
    x"ffff000000000000000b0000000000291efff5c91eff",
    x"ffff000000000000001d0000000000291efff5c913ff",
    x"ffff00000000000000150000000000291efff5c908ff",
    x"ffff00000000000000100000000000291efff5c8feff",
    x"ffff00000000000000170000000000291efff5c8f3ff",
    x"ffff00000000000000100000000000291ffff5c8e8ff",
    x"ffff00000000000000080000000000291efff5c8deff",
    x"ffff00000000000000160000000000291ffff5c8d3ff",
    x"ffff000000000000001f0000000000291ffff5c8c8ff",
    x"ffff000000000000001f0000000000291ffff5c8beff",
    x"ffff00000000000000180000000000291ffff5c8b3ff",
    x"ffff000000000000001a00000000002920fff5c8a9ff",
    x"ffff000000000000001b0000000000291ffff5c89eff",
    x"ffff000000000000001300000000002920fff5c893ff",
    x"ffff000000000000000300000000002920fff5c889ff",
    x"ffff000000000000001e00000000002920fff5c87eff",
    x"ffff000000000000001100000000002921fff5c873ff",
    x"ffff000000000000001700000000002920fff5c869ff",
    x"ffff000000000000001200000000002921fff5c85eff",
    x"ffff000000000000000100000000002923fff5c853ff",
    x"ffff000000000000001100000000002921fff5c849ff",
    x"ffff000000000000001100000000002921fff5c83eff",
    x"ffff000000000000001800000000002922fff5c833ff",
    x"ffff000000000000000e00000000002921fff5c829ff",
    x"ffff000000000000000400000000002922fff5c81eff",
    x"ffff000000000000000700000000002922fff5c814ff",
    x"ffff000000000000001b00000000002922fff5c809ff",
    x"ffff000000000000000200000000002922fff5c7feff",
    x"ffff000000000000000000000000002922fff5c7f4ff",
    x"ffff000000000000001b00000000002922fff5c7e9ff",
    x"ffff000000000000000a00000000002923fff5c7deff",
    x"ffff000000000000001500000000002923fff5c7d4ff",
    x"ffff000000000000000200000000002923fff5c7c9ff",
    x"ffff000000000000001d00000000002923fff5c7beff",
    x"ffff000000000000001400000000002923fff5c7b4ff",
    x"ffff000000000000001f00000000002924fff5c7a9ff",
    x"ffff000000000000001f00000000002923fff5c79eff",
    x"ffff000000000000001f00000000002924fff5c794ff",
    x"ffff000000000000001100000000002924fff5c789ff",
    x"ffff000000000000001a00000000002924fff5c77fff",
    x"ffff000000000000000200000000002924fff5c774ff",
    x"ffff000000000000001100000000002925fff5c769ff",
    x"ffff000000000000000600000000002925fff5c75fff",
    x"ffff000000000000000000000000002924fff5c754ff",
    x"ffff000000000000000000000000002925fff5c749ff",
    x"ffff000000000000000000000000002926fff5c73fff",
    x"ffff000000000000000900000000002925fff5c734ff",
    x"ffff000000000000000a00000000002925fff5c729ff",
    x"ffff000000000000001100000000002926fff5c71fff",
    x"ffff000000000000000500000000002926fff5c714ff",
    x"ffff000000000000000000000000002926fff5c709ff",
    x"ffff000000000000001e00000000002926fff5c6ffff",
    x"ffff000000000000000400000000002926fff5c6f4ff",
    x"ffff000000000000001c00000000002927fff5c6eaff",
    x"ffff000000000000001100000000002926fff5c6dfff",
    x"ffff000000000000000200000000002927fff5c6d4ff",
    x"ffff000000000000000000000000002927fff5c6caff",
    x"ffff000000000000001000000000002927fff5c6bfff",
    x"ffff000000000000000400000000002928fff5c6b4ff",
    x"ffff000000000000000000000000002927fff5c6aaff",
    x"ffff000000000000000000000000002928fff5c69fff",
    x"ffff000000000000000000000000002927fff5c694ff",
    x"ffff000000000000000000000000002928fff5c68aff",
    x"ffff000000000000000000000000002929fff5c67fff",
    x"ffff000000000000000000000000002928fff5c674ff",
    x"ffff000000000000000000000000002928fff5c66aff",
    x"ffff000000000000000000000000002929fff5c65fff",
    x"ffff000000000000000000000000002929fff5c655ff",
    x"ffff000000000000000000000000002929fff5c64aff",
    x"ffff000000000000000000000000002929fff5c63fff",
    x"ffff000000000000000000000000002929fff5c635ff",
    x"ffff00000000000000000000000000292afff5c62aff",
    x"ffff000000000000000000000000002929fff5c61fff",
    x"ffff00000000000000000000000000292afff5c615ff",
    x"ffff00000000000000000000000000292afff5c60aff",
    x"ffff00000000000000000000000000292afff5c5ffff",
    x"ffff00000000000000000000000000292bfff5c5f5ff",
    x"ffff00000000000000000000000000292afff5c5eaff",
    x"ffff00000000000000000000000000292bfff5c5dfff",
    x"ffff00000000000000000000000000292bfff5c5d5ff",
    x"ffff000000000000000e0000000000292bfff5c5caff",
    x"ffff00000000000000010000000000292bfff5c5c0ff",
    x"ffff000000000000001b0000000000292bfff5c5b5ff",
    x"ffff00000000000000050000000000292cfff5c5aaff",
    x"ffff00000000000000190000000000292bfff5c5a0ff",
    x"ffff000000000000001f0000000000292cfff5c595ff",
    x"ffff000000000000001f0000000000292cfff5c58aff",
    x"ffff000000000000001f0000000000292cfff5c580ff",
    x"ffff000000000000001e0000000000292dfff5c575ff",
    x"ffff000000000000001f0000000000292cfff5c56aff",
    x"ffff00000000000000070000000000292dfff5c560ff",
    x"ffff00000000000000000000000000292dfff5c555ff",
    x"ffff00000000000000000000000000292dfff5c54aff",
    x"ffff00000000000000030000000000292dfff5c540ff",
    x"ffff000000000000001d0000000000292dfff5c535ff",
    x"ffff00000000000000080000000000292efff5c52aff",
    x"ffff000000000000001e0000000000292dfff5c520ff",
    x"ffff000000000000000a0000000000292efff5c515ff",
    x"ffff00000000000000000000000000292efff5c50bff",
    x"ffff00000000000000140000000000292efff5c500ff",
    x"ffff00000000000000010000000000292ffff5c4f5ff",
    x"ffff00000000000000110000000000292efff5c4ebff",
    x"ffff00000000000000060000000000292ffff5c4e0ff",
    x"ffff00000000000000000000000000292ffff5c4d5ff",
    x"ffff00000000000000000000000000292ffff5c4cbff",
    x"ffff00000000000000000000000000292ffff5c4c0ff",
    x"ffff00000000000000090000000000292ffff5c4b5ff",
    x"ffff000000000000000a00000000002930fff5c4abff",
    x"ffff00000000000000110000000000292ffff5c4a0ff",
    x"ffff000000000000000500000000002930fff5c495ff",
    x"ffff000000000000000200000000002930fff5c48bff",
    x"ffff000000000000000500000000002930fff5c480ff",
    x"ffff000000000000000600000000002931fff5c475ff",
    x"ffff000000000000001a00000000002930fff5c46bff",
    x"ffff000000000000000600000000002931fff5c460ff",
    x"ffff000000000000001000000000002931fff5c456ff",
    x"ffff000000000000001100000000002931fff5c44bff",
    x"ffff000000000000001900000000002931fff5c440ff",
    x"ffff000000000000000200000000002931fff5c436ff",
    x"ffff000000000000000c00000000002932fff5c42bff",
    x"ffff000000000000001400000000002932fff5c420ff",
    x"ffff000000000000001e00000000002932fff5c416ff",
    x"ffff000000000000001800000000002932fff5c40bff",
    x"ffff000000000000001600000000002932fff5c400ff",
    x"ffff000000000000000d00000000002932fff5c3f6ff",
    x"ffff000000000000000200000000002933fff5c3ebff",
    x"ffff000000000000000200000000002932fff5c3e0ff",
    x"ffff000000000000000300000000002933fff5c3d6ff",
    x"ffff000000000000001900000000002933fff5c3cbff",
    x"ffff000000000000000600000000002933fff5c3c1ff",
    x"ffff000000000000001b00000000002934fff5c3b6ff",
    x"ffff000000000000001f00000000002933fff5c3abff",
    x"ffff000000000000000d00000000002934fff5c3a1ff",
    x"ffff000000000000001000000000002934fff5c396ff",
    x"ffff000000000000001e00000000002934fff5c38bff",
    x"ffff000000000000001300000000002934fff5c381ff",
    x"ffff000000000000000500000000002934fff5c376ff",
    x"ffff000000000000000000000000002935fff5c36bff",
    x"ffff000000000000000400000000002935fff5c361ff",
    x"ffff000000000000001b00000000002935fff5c356ff",
    x"ffff000000000000001500000000002935fff5c34bff",
    x"ffff000000000000000700000000002935fff5c341ff",
    x"ffff000000000000001600000000002935fff5c336ff",
    x"ffff000000000000000f00000000002936fff5c32bff",
    x"ffff000000000000000100000000002935fff5c321ff",
    x"ffff000000000000001800000000002936fff5c316ff",
    x"ffff000000000000001400000000002936fff5c30cff",
    x"ffff000000000000000700000000002937fff5c301ff",
    x"ffff000000000000000700000000002936fff5c2f6ff",
    x"ffff000000000000001000000000002936fff5c2ecff",
    x"ffff000000000000000300000000002937fff5c2e1ff",
    x"ffff000000000000001200000000002937fff5c2d6ff",
    x"ffff000000000000001f00000000002937fff5c2ccff",
    x"ffff000000000000000100000000002937fff5c2c1ff",
    x"ffff000000000000000700000000002938fff5c2b6ff",
    x"ffff000000000000001c00000000002937fff5c2acff",
    x"ffff000000000000001700000000002938fff5c2a1ff",
    x"ffff000000000000000400000000002938fff5c296ff",
    x"ffff000000000000000000000000002938fff5c28cff",
    x"ffff000000000000000c00000000002938fff5c281ff",
    x"ffff000000000000000000000000002938fff5c276ff",
    x"ffff000000000000001100000000002939fff5c26cff",
    x"ffff000000000000000600000000002939fff5c261ff",
    x"ffff000000000000000000000000002939fff5c256ff",
    x"ffff000000000000000000000000002939fff5c24cff",
    x"ffff000000000000000000000000002939fff5c241ff",
    x"ffff000000000000000900000000002939fff5c236ff",
    x"ffff000000000000000a0000000000293afff5c22cff",
    x"ffff00000000000000110000000000293afff5c221ff",
    x"ffff000000000000000500000000002939fff5c217ff",
    x"ffff00000000000000010000000000293bfff5c20cff",
    x"ffff000000000000001f0000000000293afff5c201ff",
    x"ffff00000000000000070000000000293dfff5c1f7ff",
    x"ffff000000000000001f0000000000293bfff5c1ecff",
    x"ffff000000000000001f0000000000293afff5c1e1ff",
    x"ffff00000000000000020000000000293bfff5c1d7ff",
    x"ffff00000000000000000000000000293bfff5c1ccff",
    x"ffff00000000000000120000000000293cfff5c1c1ff",
    x"ffff00000000000000100000000000293bfff5c1b7ff",
    x"ffff00000000000000180000000000293cfff5c1acff",
    x"ffff000000000000001e0000000000293bfff5c1a1ff",
    x"ffff00000000000000030000000000293cfff5c197ff",
    x"ffff000000000000001f0000000000293cfff5c18cff",
    x"ffff000000000000000d0000000000293dfff5c181ff",
    x"ffff00000000000000190000000000293cfff5c177ff",
    x"ffff00000000000000000000000000293dfff5c16cff",
    x"ffff00000000000000000000000000293cfff5c161ff",
    x"ffff00000000000000020000000000293dfff5c157ff",
    x"ffff00000000000000160000000000293dfff5c14cff",
    x"ffff00000000000000110000000000293efff5c142ff",
    x"ffff000000000000000a0000000000293dfff5c137ff",
    x"ffff000000000000001e0000000000293efff5c12cff",
    x"ffff000000000000001c0000000000293dfff5c122ff",
    x"ffff000000000000001e0000000000293efff5c117ff",
    x"ffff00000000000000040000000000293efff5c10cff",
    x"ffff00000000000000050000000000293ffff5c102ff",
    x"ffff00000000000000130000000000293efff5c0f7ff",
    x"ffff000000000000001b0000000000293efff5c0ecff",
    x"ffff00000000000000050000000000293ffff5c0e2ff",
    x"ffff000000000000000f0000000000293ffff5c0d7ff",
    x"ffff00000000000000060000000000293ffff5c0ccff",
    x"ffff000000000000000b00000000002940fff5c0c2ff",
    x"ffff00000000000000090000000000293ffff5c0b7ff",
    x"ffff000000000000001100000000002940fff5c0acff",
    x"ffff00000000000000030000000000293ffff5c0a2ff",
    x"ffff000000000000001800000000002940fff5c097ff",
    x"ffff000000000000000200000000002940fff5c08cff",
    x"ffff000000000000000900000000002941fff5c082ff",
    x"ffff000000000000001800000000002940fff5c077ff",
    x"ffff000000000000000000000000002941fff5c06cff",
    x"ffff000000000000001000000000002940fff5c062ff",
    x"ffff000000000000001600000000002941fff5c057ff",
    x"ffff000000000000001400000000002941fff5c04dff",
    x"ffff000000000000000200000000002942fff5c042ff",
    x"ffff000000000000000100000000002941fff5c037ff",
    x"ffff000000000000001a00000000002942fff5c02dff",
    x"ffff000000000000000600000000002941fff5c022ff",
    x"ffff000000000000001400000000002942fff5c017ff",
    x"ffff000000000000001c00000000002942fff5c00dff",
    x"ffff000000000000001900000000002943fff5c002ff",
    x"ffff000000000000000100000000002942fff5bff7ff",
    x"ffff000000000000001100000000002943fff5bfedff",
    x"ffff000000000000000600000000002943fff5bfe2ff",
    x"ffff000000000000000000000000002942fff5bfd7ff",
    x"ffff000000000000000000000000002944fff5bfcdff",
    x"ffff000000000000000000000000002943fff5bfc2ff",
    x"ffff000000000000000900000000002943fff5bfb7ff",
    x"ffff000000000000000a00000000002944fff5bfadff",
    x"ffff000000000000001100000000002944fff5bfa2ff",
    x"ffff000000000000000500000000002944fff5bf97ff",
    x"ffff000000000000001300000000002944fff5bf8dff",
    x"ffff000000000000001400000000002944fff5bf82ff",
    x"ffff000000000000000300000000002944fff5bf77ff",
    x"ffff000000000000001d00000000002945fff5bf6dff",
    x"ffff000000000000000400000000002945fff5bf62ff",
    x"ffff000000000000000000000000002945fff5bf58ff",
    x"ffff000000000000000000000000002945fff5bf4dff",
    x"ffff000000000000001000000000002945fff5bf42ff",
    x"ffff000000000000001e00000000002946fff5bf38ff",
    x"ffff000000000000001f00000000002945fff5bf2dff",
    x"ffff000000000000001f00000000002946fff5bf22ff",
    x"ffff000000000000001f00000000002946fff5bf18ff",
    x"ffff000000000000001f00000000002946fff5bf0dff",
    x"ffff000000000000001f00000000002946fff5bf02ff",
    x"ffff000000000000001f00000000002947fff5bef8ff",
    x"ffff000000000000001f00000000002946fff5beedff",
    x"ffff000000000000001f00000000002947fff5bee2ff",
    x"ffff000000000000001f00000000002947fff5bed8ff",
    x"ffff000000000000001f00000000002947fff5becdff",
    x"ffff000000000000001f00000000002948fff5bec2ff",
    x"ffff000000000000001f00000000002947fff5beb8ff",
    x"ffff000000000000001f00000000002948fff5beadff",
    x"ffff000000000000001f00000000002948fff5bea2ff",
    x"ffff000000000000001f00000000002948fff5be98ff",
    x"ffff000000000000001f00000000002948fff5be8dff",
    x"ffff000000000000001f00000000002948fff5be82ff",
    x"ffff000000000000001f00000000002948fff5be78ff",
    x"ffff000000000000001f00000000002949fff5be6dff",
    x"ffff000000000000001f00000000002949fff5be62ff",
    x"ffff000000000000001f00000000002949fff5be58ff",
    x"ffff000000000000001f00000000002949fff5be4dff",
    x"ffff000000000000001f00000000002949fff5be43ff",
    x"ffff000000000000001f0000000000294afff5be38ff",
    x"ffff000000000000001f00000000002949fff5be2dff",
    x"ffff000000000000001f0000000000294afff5be23ff",
    x"ffff000000000000001f0000000000294afff5be18ff",
    x"ffff000000000000001f0000000000294afff5be0dff",
    x"ffff000000000000001f0000000000294bfff5be03ff",
    x"ffff000000000000001f0000000000294afff5bdf8ff",
    x"ffff000000000000001f0000000000294bfff5bdedff",
    x"ffff000000000000001f0000000000294afff5bde3ff",
    x"ffff000000000000001f0000000000294bfff5bdd8ff",
    x"ffff000000000000001f0000000000294cfff5bdcdff",
    x"ffff000000000000001f0000000000294bfff5bdc3ff",
    x"ffff000000000000001f0000000000294bfff5bdb8ff",
    x"ffff000000000000001f0000000000294cfff5bdadff",
    x"ffff000000000000001f0000000000294cfff5bda3ff",
    x"ffff000000000000001f0000000000294cfff5bd98ff",
    x"ffff000000000000001f0000000000294cfff5bd8dff",
    x"ffff00000000000000170000000000294cfff5bd83ff",
    x"ffff00000000000000060000000000294dfff5bd78ff",
    x"ffff00000000000000110000000000294cfff5bd6dff",
    x"ffff00000000000000060000000000294dfff5bd63ff",
    x"ffff00000000000000000000000000294dfff5bd58ff",
    x"ffff00000000000000000000000000294dfff5bd4dff",
    x"ffff00000000000000000000000000294efff5bd43ff",
    x"ffff00000000000000090000000000294dfff5bd38ff",
    x"ffff000000000000000a0000000000294efff5bd2dff",
    x"ffff00000000000000110000000000294efff5bd23ff",
    x"ffff00000000000000150000000000294efff5bd18ff",
    x"ffff00000000000000100000000000294efff5bd0eff",
    x"ffff00000000000000060000000000294efff5bd03ff",
    x"ffff00000000000000040000000000294ffff5bcf8ff",
    x"ffff00000000000000120000000000294efff5bceeff",
    x"ffff00000000000000050000000000294ffff5bce3ff",
    x"ffff000000000000001f0000000000294ffff5bcd8ff",
    x"ffff00000000000000110000000000294ffff5bcceff",
    x"ffff000000000000001c00000000002950fff5bcc3ff",
    x"ffff00000000000000000000000000294ffff5bcb8ff",
    x"ffff000000000000000000000000002950fff5bcaeff",
    x"ffff000000000000000400000000002950fff5bca3ff",
    x"ffff000000000000000700000000002950fff5bc98ff",
    x"ffff000000000000000a00000000002950fff5bc8eff",
    x"ffff000000000000001e00000000002950fff5bc83ff",
    x"ffff000000000000001b00000000002951fff5bc78ff",
    x"ffff000000000000001000000000002950fff5bc6eff",
    x"ffff000000000000000800000000002951fff5bc63ff",
    x"ffff000000000000000b00000000002951fff5bc58ff",
    x"ffff000000000000001f00000000002951fff5bc4eff",
    x"ffff000000000000001f00000000002952fff5bc43ff",
    x"ffff000000000000001c00000000002951fff5bc38ff",
    x"ffff000000000000001a00000000002952fff5bc2eff",
    x"ffff000000000000001b00000000002952fff5bc23ff",
    x"ffff000000000000001300000000002952fff5bc18ff",
    x"ffff000000000000001a00000000002952fff5bc0eff",
    x"ffff000000000000000400000000002952fff5bc03ff",
    x"ffff000000000000000900000000002953fff5bbf8ff",
    x"ffff000000000000001500000000002953fff5bbeeff",
    x"ffff000000000000001500000000002952fff5bbe3ff",
    x"ffff000000000000000400000000002954fff5bbd8ff",
    x"ffff000000000000000900000000002953fff5bbceff",
    x"ffff000000000000000400000000002953fff5bbc3ff",
    x"ffff000000000000001000000000002954fff5bbb8ff",
    x"ffff000000000000000100000000002953fff5bbaeff",
    x"ffff000000000000000d00000000002954fff5bba3ff",
    x"ffff000000000000000b00000000002957fff5bb98ff",
    x"ffff000000000000000d00000000002954fff5bb8eff",
    x"ffff000000000000001f00000000002955fff5bb83ff",
    x"ffff000000000000001b00000000002954fff5bb78ff",
    x"ffff000000000000001500000000002955fff5bb6eff",
    x"ffff000000000000001100000000002955fff5bb63ff",
    x"ffff000000000000001700000000002955fff5bb59ff",
    x"ffff000000000000000600000000002955fff5bb4eff",
    x"ffff000000000000000600000000002955fff5bb43ff",
    x"ffff000000000000001c00000000002956fff5bb39ff",
    x"ffff000000000000000d00000000002956fff5bb2eff",
    x"ffff000000000000001c00000000002955fff5bb23ff",
    x"ffff000000000000001f00000000002956fff5bb19ff",
    x"ffff000000000000001700000000002957fff5bb0eff",
    x"ffff000000000000001800000000002956fff5bb03ff",
    x"ffff000000000000000200000000002957fff5baf9ff",
    x"ffff000000000000001100000000002956fff5baeeff",
    x"ffff000000000000000600000000002957fff5bae3ff",
    x"ffff000000000000000000000000002957fff5bad9ff",
    x"ffff000000000000000000000000002958fff5baceff",
    x"ffff000000000000000000000000002957fff5bac3ff",
    x"ffff000000000000000900000000002957fff5bab9ff",
    x"ffff000000000000000a00000000002958fff5baaeff",
    x"ffff000000000000001100000000002958fff5baa3ff",
    x"ffff000000000000001500000000002958fff5ba99ff",
    x"ffff000000000000000200000000002958fff5ba8eff",
    x"ffff000000000000001a00000000002959fff5ba83ff",
    x"ffff000000000000000300000000002958fff5ba79ff",
    x"ffff000000000000001c00000000002959fff5ba6eff",
    x"ffff000000000000001100000000002959fff5ba63ff",
    x"ffff000000000000000200000000002959fff5ba59ff",
    x"ffff000000000000000000000000002959fff5ba4eff",
    x"ffff000000000000001000000000002959fff5ba43ff",
    x"ffff00000000000000040000000000295afff5ba39ff",
    x"ffff00000000000000000000000000295afff5ba2eff",
    x"ffff00000000000000000000000000295afff5ba23ff",
    x"ffff00000000000000000000000000295afff5ba19ff",
    x"ffff00000000000000000000000000295afff5ba0eff",
    x"ffff00000000000000000000000000295afff5ba03ff",
    x"ffff00000000000000000000000000295bfff5b9f9ff",
    x"ffff00000000000000000000000000295bfff5b9eeff",
    x"ffff00000000000000000000000000295bfff5b9e3ff",
    x"ffff00000000000000000000000000295bfff5b9d9ff",
    x"ffff00000000000000000000000000295bfff5b9ceff",
    x"ffff00000000000000000000000000295bfff5b9c3ff",
    x"ffff00000000000000000000000000295cfff5b9b9ff",
    x"ffff00000000000000000000000000295cfff5b9aeff",
    x"ffff00000000000000000000000000295cfff5b9a3ff",
    x"ffff00000000000000000000000000295cfff5b999ff",
    x"ffff00000000000000000000000000295cfff5b98eff",
    x"ffff00000000000000000000000000295cfff5b983ff",
    x"ffff00000000000000000000000000295dfff5b979ff",
    x"ffff00000000000000000000000000295dfff5b96eff",
    x"ffff00000000000000000000000000295cfff5b963ff",
    x"ffff00000000000000000000000000295efff5b959ff",
    x"ffff000000000000000e0000000000295dfff5b94eff",
    x"ffff00000000000000010000000000295dfff5b943ff",
    x"ffff000000000000001b0000000000295efff5b939ff",
    x"ffff00000000000000050000000000295efff5b92eff",
    x"ffff00000000000000190000000000295dfff5b923ff",
    x"ffff000000000000001f0000000000295ffff5b919ff",
    x"ffff000000000000001f0000000000295efff5b90eff",
    x"ffff000000000000001f0000000000295efff5b903ff",
    x"ffff000000000000001e0000000000295ffff5b8f9ff",
    x"ffff000000000000001f0000000000295ffff5b8eeff",
    x"ffff00000000000000070000000000295efff5b8e4ff",
    x"ffff000000000000000000000000002960fff5b8d9ff",
    x"ffff00000000000000000000000000295ffff5b8ceff",
    x"ffff00000000000000030000000000295ffff5b8c4ff",
    x"ffff000000000000001d00000000002960fff5b8b9ff",
    x"ffff000000000000000800000000002960fff5b8aeff",
    x"ffff000000000000001e0000000000295ffff5b8a4ff",
    x"ffff000000000000000a00000000002961fff5b899ff",
    x"ffff000000000000000000000000002960fff5b88eff",
    x"ffff000000000000001400000000002960fff5b884ff",
    x"ffff000000000000000100000000002961fff5b879ff",
    x"ffff000000000000001100000000002961fff5b86eff",
    x"ffff000000000000000600000000002961fff5b864ff",
    x"ffff000000000000000000000000002961fff5b859ff",
    x"ffff000000000000000000000000002961fff5b84eff",
    x"ffff000000000000000000000000002961fff5b844ff",
    x"ffff000000000000000900000000002962fff5b839ff",
    x"ffff000000000000000a00000000002962fff5b82eff",
    x"ffff000000000000001100000000002962fff5b824ff",
    x"ffff000000000000001500000000002962fff5b819ff",
    x"ffff000000000000000100000000002962fff5b80eff",
    x"ffff000000000000001d00000000002963fff5b804ff",
    x"ffff000000000000000200000000002962fff5b7f9ff",
    x"ffff000000000000001a00000000002963fff5b7eeff",
    x"ffff000000000000000600000000002963fff5b7e4ff",
    x"ffff000000000000001000000000002963fff5b7d9ff",
    x"ffff000000000000001100000000002963fff5b7ceff",
    x"ffff000000000000001900000000002964fff5b7c4ff",
    x"ffff000000000000000200000000002963fff5b7b9ff",
    x"ffff000000000000000c00000000002964fff5b7aeff",
    x"ffff000000000000001400000000002964fff5b7a4ff",
    x"ffff000000000000001e00000000002964fff5b799ff",
    x"ffff000000000000001800000000002965fff5b78eff",
    x"ffff000000000000001600000000002964fff5b784ff",
    x"ffff000000000000000d00000000002965fff5b779ff",
    x"ffff000000000000000200000000002964fff5b76eff",
    x"ffff000000000000000200000000002965fff5b764ff",
    x"ffff000000000000000300000000002965fff5b759ff",
    x"ffff000000000000001900000000002966fff5b74eff",
    x"ffff000000000000000600000000002965fff5b744ff",
    x"ffff000000000000001b00000000002966fff5b739ff",
    x"ffff000000000000001f00000000002966fff5b72eff",
    x"ffff000000000000000d00000000002966fff5b724ff",
    x"ffff000000000000001000000000002966fff5b719ff",
    x"ffff000000000000001e00000000002966fff5b70eff",
    x"ffff000000000000001300000000002967fff5b704ff",
    x"ffff000000000000000500000000002966fff5b6f9ff",
    x"ffff000000000000000000000000002967fff5b6eeff",
    x"ffff000000000000000400000000002967fff5b6e4ff",
    x"ffff000000000000001b00000000002967fff5b6d9ff",
    x"ffff000000000000001500000000002968fff5b6ceff",
    x"ffff000000000000000700000000002967fff5b6c4ff",
    x"ffff000000000000001600000000002968fff5b6b9ff",
    x"ffff000000000000000f00000000002967fff5b6aeff",
    x"ffff000000000000000100000000002968fff5b6a4ff",
    x"ffff000000000000001800000000002969fff5b699ff",
    x"ffff000000000000001400000000002968fff5b68eff",
    x"ffff000000000000000700000000002968fff5b684ff",
    x"ffff000000000000000700000000002969fff5b679ff",
    x"ffff000000000000001000000000002969fff5b66eff",
    x"ffff000000000000000300000000002969fff5b664ff",
    x"ffff000000000000001200000000002969fff5b659ff",
    x"ffff000000000000001f00000000002969fff5b64eff",
    x"ffff00000000000000010000000000296afff5b644ff",
    x"ffff000000000000000700000000002969fff5b639ff",
    x"ffff000000000000001c0000000000296afff5b62eff",
    x"ffff00000000000000170000000000296afff5b624ff",
    x"ffff00000000000000040000000000296afff5b619ff",
    x"ffff00000000000000000000000000296bfff5b60eff",
    x"ffff000000000000000c0000000000296afff5b604ff",
    x"ffff00000000000000000000000000296bfff5b5f9ff",
    x"ffff00000000000000110000000000296bfff5b5eeff",
    x"ffff00000000000000060000000000296bfff5b5e4ff",
    x"ffff00000000000000000000000000296bfff5b5d9ff",
    x"ffff00000000000000000000000000296bfff5b5ceff",
    x"ffff00000000000000000000000000296cfff5b5c4ff",
    x"ffff00000000000000090000000000296bfff5b5b9ff",
    x"ffff000000000000000a0000000000296cfff5b5aeff",
    x"ffff00000000000000110000000000296cfff5b5a4ff",
    x"ffff00000000000000150000000000296cfff5b599ff",
    x"ffff00000000000000030000000000296dfff5b58eff",
    x"ffff000000000000001b0000000000296cfff5b584ff",
    x"ffff00000000000000000000000000296dfff5b579ff",
    x"ffff000000000000001f0000000000296dfff5b56eff",
    x"ffff000000000000001f0000000000296dfff5b564ff",
    x"ffff00000000000000020000000000296dfff5b559ff",
    x"ffff00000000000000000000000000296dfff5b54eff",
    x"ffff00000000000000120000000000296efff5b544ff",
    x"ffff000000000000001000000000002970fff5b539ff",
    x"ffff00000000000000180000000000296efff5b52eff",
    x"ffff000000000000001e0000000000296efff5b524ff",
    x"ffff00000000000000030000000000296ffff5b519ff",
    x"ffff000000000000001f0000000000296efff5b50eff",
    x"ffff000000000000000d0000000000296efff5b504ff",
    x"ffff00000000000000190000000000296ffff5b4f9ff",
    x"ffff00000000000000000000000000296ffff5b4eeff",
    x"ffff00000000000000000000000000296ffff5b4e4ff",
    x"ffff00000000000000020000000000296ffff5b4d9ff",
    x"ffff00000000000000160000000000296ffff5b4ceff",
    x"ffff000000000000001100000000002970fff5b4c4ff",
    x"ffff000000000000000a00000000002970fff5b4b9ff",
    x"ffff000000000000001e00000000002970fff5b4aeff",
    x"ffff000000000000001c00000000002970fff5b4a4ff",
    x"ffff000000000000001e00000000002970fff5b499ff",
    x"ffff000000000000000400000000002970fff5b48eff",
    x"ffff000000000000000500000000002971fff5b484ff",
    x"ffff000000000000001300000000002970fff5b479ff",
    x"ffff000000000000001b00000000002971fff5b46eff",
    x"ffff000000000000000500000000002971fff5b464ff",
    x"ffff000000000000000f00000000002972fff5b459ff",
    x"ffff000000000000000600000000002971fff5b44eff",
    x"ffff000000000000000b00000000002971fff5b444ff",
    x"ffff000000000000000900000000002972fff5b439ff",
    x"ffff000000000000001100000000002972fff5b42eff",
    x"ffff000000000000000300000000002972fff5b424ff",
    x"ffff000000000000001800000000002972fff5b419ff",
    x"ffff000000000000000200000000002973fff5b40eff",
    x"ffff000000000000000900000000002972fff5b404ff",
    x"ffff000000000000001800000000002973fff5b3f9ff",
    x"ffff000000000000000000000000002973fff5b3eeff",
    x"ffff000000000000001000000000002973fff5b3e4ff",
    x"ffff000000000000001600000000002973fff5b3d9ff",
    x"ffff000000000000001400000000002973fff5b3ceff",
    x"ffff000000000000000200000000002974fff5b3c4ff",
    x"ffff000000000000000100000000002974fff5b3b9ff",
    x"ffff000000000000001a00000000002974fff5b3aeff",
    x"ffff000000000000000600000000002974fff5b3a4ff",
    x"ffff000000000000001400000000002974fff5b399ff",
    x"ffff000000000000001c00000000002974fff5b38eff",
    x"ffff000000000000001900000000002975fff5b384ff",
    x"ffff000000000000000100000000002975fff5b379ff",
    x"ffff000000000000001100000000002974fff5b36eff",
    x"ffff000000000000000600000000002975fff5b364ff",
    x"ffff000000000000000000000000002976fff5b359ff",
    x"ffff000000000000000000000000002975fff5b34eff",
    x"ffff000000000000000000000000002976fff5b344ff",
    x"ffff000000000000000900000000002975fff5b339ff",
    x"ffff000000000000000a00000000002976fff5b32eff",
    x"ffff000000000000001100000000002976fff5b324ff",
    x"ffff000000000000000d00000000002977fff5b319ff",
    x"ffff000000000000001000000000002976fff5b30eff",
    x"ffff000000000000000800000000002977fff5b303ff",
    x"ffff000000000000000300000000002976fff5b2f9ff",
    x"ffff000000000000001d00000000002977fff5b2eeff",
    x"ffff000000000000000400000000002977fff5b2e3ff",
    x"ffff000000000000000000000000002978fff5b2d9ff",
    x"ffff000000000000000000000000002977fff5b2ceff",
    x"ffff000000000000001000000000002978fff5b2c3ff",
    x"ffff000000000000001e00000000002977fff5b2b9ff",
    x"ffff000000000000001f00000000002978fff5b2aeff",
    x"ffff000000000000001f00000000002978fff5b2a3ff",
    x"ffff000000000000001f00000000002979fff5b299ff",
    x"ffff000000000000001f00000000002978fff5b28eff",
    x"ffff000000000000001f00000000002979fff5b283ff",
    x"ffff000000000000001f00000000002978fff5b279ff",
    x"ffff000000000000001f00000000002979fff5b26eff",
    x"ffff000000000000001f00000000002979fff5b263ff",
    x"ffff000000000000001f0000000000297afff5b259ff",
    x"ffff000000000000001f00000000002979fff5b24eff",
    x"ffff000000000000001f0000000000297afff5b243ff",
    x"ffff000000000000001f00000000002979fff5b239ff",
    x"ffff000000000000001f0000000000297afff5b22eff",
    x"ffff000000000000001f0000000000297afff5b223ff",
    x"ffff000000000000001f0000000000297bfff5b219ff",
    x"ffff000000000000001f0000000000297afff5b20eff",
    x"ffff000000000000001f0000000000297bfff5b203ff",
    x"ffff000000000000001f0000000000297afff5b1f9ff",
    x"ffff000000000000001f0000000000297bfff5b1eeff",
    x"ffff000000000000001f0000000000297cfff5b1e3ff",
    x"ffff000000000000001f0000000000297bfff5b1d9ff",
    x"ffff000000000000001f0000000000297bfff5b1ceff",
    x"ffff000000000000001f0000000000297cfff5b1c3ff",
    x"ffff000000000000001f0000000000297cfff5b1b9ff",
    x"ffff000000000000001f0000000000297cfff5b1aeff",
    x"ffff000000000000001f0000000000297cfff5b1a3ff",
    x"ffff000000000000001f0000000000297cfff5b199ff",
    x"ffff000000000000001f0000000000297cfff5b18eff",
    x"ffff000000000000001f0000000000297dfff5b183ff",
    x"ffff000000000000001f0000000000297dfff5b179ff",
    x"ffff000000000000001f0000000000297dfff5b16eff",
    x"ffff000000000000001f0000000000297dfff5b163ff",
    x"ffff000000000000001f0000000000297dfff5b159ff",
    x"ffff000000000000001f0000000000297efff5b14eff",
    x"ffff000000000000001f0000000000297dfff5b143ff",
    x"ffff000000000000001f0000000000297efff5b139ff",
    x"ffff000000000000001f0000000000297efff5b12eff",
    x"ffff000000000000001f0000000000297efff5b123ff",
    x"ffff000000000000001f0000000000297efff5b119ff",
    x"ffff000000000000001f0000000000297ffff5b10eff",
    x"ffff00000000000000170000000000297efff5b103ff",
    x"ffff00000000000000060000000000297ffff5b0f9ff",
    x"ffff00000000000000110000000000297ffff5b0eeff",
    x"ffff00000000000000060000000000297ffff5b0e3ff",
    x"ffff000000000000000000000000002980fff5b0d8ff",
    x"ffff00000000000000000000000000297ffff5b0ceff",
    x"ffff000000000000000000000000002980fff5b0c3ff",
    x"ffff000000000000000900000000002980fff5b0b8ff",
    x"ffff000000000000000a00000000002980fff5b0aeff",
    x"ffff000000000000001100000000002980fff5b0a3ff",
    x"ffff000000000000000d00000000002980fff5b098ff",
    x"ffff000000000000001200000000002980fff5b08eff",
    x"ffff000000000000000e00000000002981fff5b083ff",
    x"ffff000000000000000100000000002981fff5b078ff",
    x"ffff000000000000000a00000000002981fff5b06eff",
    x"ffff000000000000000700000000002981fff5b063ff",
    x"ffff000000000000001e00000000002981fff5b058ff",
    x"ffff000000000000000700000000002982fff5b04eff",
    x"ffff000000000000001a00000000002981fff5b043ff",
    x"ffff000000000000000e00000000002982fff5b038ff",
    x"ffff000000000000000000000000002982fff5b02eff",
    x"ffff000000000000001400000000002982fff5b023ff",
    x"ffff000000000000001800000000002983fff5b018ff",
    x"ffff000000000000000800000000002982fff5b00eff",
    x"ffff000000000000001200000000002983fff5b003ff",
    x"ffff000000000000000500000000002983fff5aff8ff",
    x"ffff000000000000000f00000000002983fff5afeeff",
    x"ffff000000000000001700000000002983fff5afe3ff",
    x"ffff000000000000000e00000000002983fff5afd8ff",
    x"ffff000000000000000000000000002984fff5afceff",
    x"ffff000000000000000000000000002983fff5afc3ff",
    x"ffff000000000000001000000000002984fff5afb8ff",
    x"ffff000000000000001a00000000002984fff5afaeff",
    x"ffff000000000000001b00000000002984fff5afa3ff",
    x"ffff000000000000001300000000002985fff5af98ff",
    x"ffff000000000000001c00000000002984fff5af8eff",
    x"ffff000000000000000a00000000002985fff5af83ff",
    x"ffff000000000000000900000000002985fff5af78ff",
    x"ffff000000000000000800000000002985fff5af6eff",
    x"ffff000000000000000c00000000002985fff5af63ff",
    x"ffff000000000000001300000000002985fff5af58ff",
    x"ffff000000000000000400000000002986fff5af4eff",
    x"ffff000000000000000b00000000002985fff5af43ff",
    x"ffff000000000000001500000000002986fff5af38ff",
    x"ffff000000000000000100000000002986fff5af2eff",
    x"ffff000000000000000900000000002986fff5af23ff",
    x"ffff000000000000000200000000002987fff5af18ff",
    x"ffff000000000000001500000000002986fff5af0dff",
    x"ffff000000000000001800000000002987fff5af03ff",
    x"ffff000000000000000500000000002987fff5aef8ff",
    x"ffff000000000000000f00000000002987fff5aeedff",
    x"ffff000000000000000f00000000002987fff5aee3ff",
    x"ffff000000000000001b00000000002987fff5aed8ff",
    x"ffff000000000000001f0000000000298bfff5aecdff",
    x"ffff000000000000001600000000002988fff5aec3ff",
    x"ffff000000000000001d00000000002987fff5aeb8ff",
    x"ffff000000000000000f00000000002989fff5aeadff",
    x"ffff000000000000001a00000000002988fff5aea3ff",
    x"ffff000000000000001f00000000002988fff5ae98ff",
    x"ffff000000000000000b00000000002989fff5ae8dff",
    x"ffff000000000000001f00000000002988fff5ae83ff",
    x"ffff000000000000000500000000002989fff5ae78ff",
    x"ffff000000000000001100000000002989fff5ae6dff",
    x"ffff000000000000000600000000002989fff5ae63ff",
    x"ffff00000000000000000000000000298afff5ae58ff",
    x"ffff000000000000000000000000002989fff5ae4dff",
    x"ffff00000000000000000000000000298afff5ae43ff",
    x"ffff00000000000000090000000000298afff5ae38ff",
    x"ffff000000000000000a0000000000298afff5ae2dff",
    x"ffff00000000000000110000000000298afff5ae23ff",
    x"ffff000000000000000d0000000000298bfff5ae18ff",
    x"ffff00000000000000010000000000298afff5ae0dff",
    x"ffff000000000000000e0000000000298bfff5ae03ff",
    x"ffff00000000000000050000000000298bfff5adf8ff",
    x"ffff000000000000001c0000000000298bfff5adedff",
    x"ffff00000000000000110000000000298bfff5ade3ff",
    x"ffff00000000000000020000000000298bfff5add8ff",
    x"ffff00000000000000000000000000298cfff5adcdff",
    x"ffff00000000000000100000000000298cfff5adc2ff",
    x"ffff00000000000000040000000000298cfff5adb8ff",
    x"ffff00000000000000000000000000298cfff5adadff",
    x"ffff00000000000000000000000000298cfff5ada2ff",
    x"ffff00000000000000000000000000298cfff5ad98ff",
    x"ffff00000000000000000000000000298dfff5ad8dff",
    x"ffff00000000000000000000000000298cfff5ad82ff",
    x"ffff00000000000000000000000000298dfff5ad78ff",
    x"ffff00000000000000000000000000298dfff5ad6dff",
    x"ffff00000000000000000000000000298efff5ad62ff",
    x"ffff00000000000000000000000000298dfff5ad58ff",
    x"ffff00000000000000000000000000298efff5ad4dff",
    x"ffff00000000000000000000000000298dfff5ad42ff",
    x"ffff00000000000000000000000000298efff5ad38ff",
    x"ffff00000000000000000000000000298efff5ad2dff",
    x"ffff00000000000000000000000000298ffff5ad22ff",
    x"ffff00000000000000000000000000298efff5ad18ff",
    x"ffff00000000000000000000000000298ffff5ad0dff",
    x"ffff00000000000000000000000000298efff5ad02ff",
    x"ffff00000000000000000000000000298ffff5acf8ff",
    x"ffff00000000000000000000000000298ffff5acedff",
    x"ffff000000000000000000000000002990fff5ace2ff",
    x"ffff00000000000000000000000000298ffff5acd8ff",
    x"ffff000000000000000e00000000002990fff5accdff",
    x"ffff00000000000000010000000000298ffff5acc2ff",
    x"ffff000000000000001b00000000002990fff5acb8ff",
    x"ffff000000000000000500000000002990fff5acadff",
    x"ffff000000000000001900000000002991fff5aca2ff",
    x"ffff000000000000001f00000000002990fff5ac97ff",
    x"ffff000000000000001f00000000002991fff5ac8dff",
    x"ffff000000000000001f00000000002990fff5ac82ff",
    x"ffff000000000000001e00000000002991fff5ac77ff",
    x"ffff000000000000001f00000000002991fff5ac6dff",
    x"ffff000000000000000700000000002992fff5ac62ff",
    x"ffff000000000000000000000000002991fff5ac57ff",
    x"ffff000000000000000000000000002992fff5ac4dff",
    x"ffff000000000000000300000000002991fff5ac42ff",
    x"ffff000000000000001d00000000002992fff5ac37ff",
    x"ffff000000000000000800000000002993fff5ac2dff",
    x"ffff000000000000001e00000000002992fff5ac22ff",
    x"ffff000000000000000a00000000002992fff5ac17ff",
    x"ffff000000000000000000000000002993fff5ac0dff",
    x"ffff000000000000001400000000002993fff5ac02ff",
    x"ffff000000000000000100000000002993fff5abf7ff",
    x"ffff000000000000001100000000002993fff5abedff",
    x"ffff000000000000000600000000002993fff5abe2ff",
    x"ffff000000000000000000000000002993fff5abd7ff",
    x"ffff000000000000000000000000002994fff5abcdff",
    x"ffff000000000000000000000000002994fff5abc2ff",
    x"ffff000000000000000900000000002994fff5abb7ff",
    x"ffff000000000000000a00000000002994fff5abacff",
    x"ffff000000000000001100000000002994fff5aba2ff",
    x"ffff000000000000000d00000000002995fff5ab97ff",
    x"ffff000000000000000300000000002994fff5ab8cff",
    x"ffff000000000000001500000000002995fff5ab82ff",
    x"ffff000000000000000700000000002995fff5ab77ff",
    x"ffff000000000000001a00000000002995fff5ab6cff",
    x"ffff000000000000000600000000002995fff5ab62ff",
    x"ffff000000000000001000000000002996fff5ab57ff",
    x"ffff000000000000001100000000002995fff5ab4cff",
    x"ffff000000000000001900000000002996fff5ab42ff",
    x"ffff000000000000000200000000002996fff5ab37ff",
    x"ffff000000000000000c00000000002996fff5ab2cff",
    x"ffff000000000000001400000000002997fff5ab22ff",
    x"ffff000000000000001e00000000002996fff5ab17ff",
    x"ffff000000000000001800000000002997fff5ab0cff",
    x"ffff000000000000001600000000002997fff5ab02ff",
    x"ffff000000000000000d00000000002997fff5aaf7ff",
    x"ffff000000000000000200000000002997fff5aaecff",
    x"ffff000000000000000200000000002997fff5aae2ff",
    x"ffff000000000000000300000000002997fff5aad7ff",
    x"ffff000000000000001900000000002998fff5aaccff",
    x"ffff000000000000000600000000002998fff5aac2ff",
    x"ffff000000000000001b00000000002998fff5aab7ff",
    x"ffff000000000000001f00000000002998fff5aaacff",
    x"ffff000000000000000d00000000002998fff5aaa1ff",
    x"ffff000000000000001000000000002999fff5aa97ff",
    x"ffff000000000000001e00000000002998fff5aa8cff",
    x"ffff000000000000001300000000002999fff5aa81ff",
    x"ffff000000000000000500000000002999fff5aa77ff",
    x"ffff000000000000000000000000002999fff5aa6cff",
    x"ffff00000000000000040000000000299afff5aa61ff",
    x"ffff000000000000001b00000000002999fff5aa57ff",
    x"ffff00000000000000150000000000299afff5aa4cff",
    x"ffff00000000000000070000000000299afff5aa41ff",
    x"ffff00000000000000160000000000299afff5aa37ff",
    x"ffff000000000000000f0000000000299afff5aa2cff",
    x"ffff00000000000000010000000000299afff5aa21ff",
    x"ffff00000000000000180000000000299bfff5aa17ff",
    x"ffff00000000000000140000000000299afff5aa0cff",
    x"ffff00000000000000070000000000299bfff5aa01ff",
    x"ffff00000000000000070000000000299bfff5a9f7ff",
    x"ffff00000000000000100000000000299bfff5a9ecff",
    x"ffff00000000000000030000000000299cfff5a9e1ff",
    x"ffff00000000000000120000000000299bfff5a9d6ff",
    x"ffff000000000000001f0000000000299cfff5a9ccff",
    x"ffff00000000000000010000000000299cfff5a9c1ff",
    x"ffff00000000000000070000000000299cfff5a9b6ff",
    x"ffff000000000000001c0000000000299cfff5a9acff",
    x"ffff00000000000000170000000000299cfff5a9a1ff",
    x"ffff00000000000000040000000000299dfff5a996ff",
    x"ffff00000000000000000000000000299dfff5a98cff",
    x"ffff000000000000000c0000000000299cfff5a981ff",
    x"ffff00000000000000000000000000299dfff5a976ff",
    x"ffff00000000000000110000000000299efff5a96cff",
    x"ffff00000000000000060000000000299dfff5a961ff",
    x"ffff00000000000000000000000000299dfff5a956ff",
    x"ffff00000000000000000000000000299efff5a94cff",
    x"ffff00000000000000000000000000299efff5a941ff",
    x"ffff00000000000000090000000000299efff5a936ff",
    x"ffff000000000000000a0000000000299efff5a92cff",
    x"ffff00000000000000110000000000299ffff5a921ff",
    x"ffff000000000000001d0000000000299efff5a916ff",
    x"ffff00000000000000000000000000299ffff5a90bff",
    x"ffff00000000000000070000000000299ffff5a901ff",
    x"ffff00000000000000000000000000299ffff5a8f6ff",
    x"ffff000000000000001f0000000000299ffff5a8ebff",
    x"ffff000000000000001f0000000000299ffff5a8e1ff",
    x"ffff0000000000000002000000000029a0fff5a8d6ff",
    x"ffff0000000000000000000000000029a0fff5a8cbff",
    x"ffff0000000000000012000000000029a0fff5a8c1ff",
    x"ffff0000000000000010000000000029a0fff5a8b6ff",
    x"ffff0000000000000018000000000029a0fff5a8abff",
    x"ffff000000000000001e000000000029a0fff5a8a1ff",
    x"ffff0000000000000003000000000029a1fff5a896ff",
    x"ffff000000000000001f000000000029a0fff5a88bff",
    x"ffff000000000000000d000000000029a1fff5a881ff",
    x"ffff0000000000000019000000000029a1fff5a876ff",
    x"ffff0000000000000000000000000029a2fff5a86bff",
    x"ffff0000000000000000000000000029a4fff5a860ff",
    x"ffff0000000000000002000000000029a2fff5a856ff",
    x"ffff0000000000000016000000000029a1fff5a84bff",
    x"ffff0000000000000011000000000029a2fff5a840ff",
    x"ffff000000000000000a000000000029a2fff5a836ff",
    x"ffff000000000000001e000000000029a2fff5a82bff",
    x"ffff000000000000001c000000000029a3fff5a820ff",
    x"ffff000000000000001e000000000029a2fff5a816ff",
    x"ffff0000000000000004000000000029a3fff5a80bff",
    x"ffff0000000000000005000000000029a3fff5a800ff",
    x"ffff0000000000000013000000000029a3fff5a7f6ff",
    x"ffff000000000000001b000000000029a3fff5a7ebff",
    x"ffff0000000000000005000000000029a4fff5a7e0ff",
    x"ffff000000000000000f000000000029a3fff5a7d6ff",
    x"ffff0000000000000006000000000029a4fff5a7cbff",
    x"ffff000000000000000b000000000029a4fff5a7c0ff",
    x"ffff0000000000000009000000000029a4fff5a7b6ff",
    x"ffff0000000000000011000000000029a4fff5a7abff",
    x"ffff0000000000000003000000000029a5fff5a7a0ff",
    x"ffff0000000000000018000000000029a4fff5a795ff",
    x"ffff0000000000000002000000000029a5fff5a78bff",
    x"ffff0000000000000009000000000029a5fff5a780ff",
    x"ffff0000000000000018000000000029a5fff5a775ff",
    x"ffff0000000000000000000000000029a5fff5a76bff",
    x"ffff0000000000000010000000000029a6fff5a760ff",
    x"ffff0000000000000016000000000029a5fff5a755ff",
    x"ffff0000000000000014000000000029a6fff5a74bff",
    x"ffff0000000000000002000000000029a6fff5a740ff",
    x"ffff0000000000000001000000000029a6fff5a735ff",
    x"ffff000000000000001a000000000029a6fff5a72bff",
    x"ffff0000000000000006000000000029a7fff5a720ff",
    x"ffff0000000000000014000000000029a6fff5a715ff",
    x"ffff000000000000001c000000000029a7fff5a70bff",
    x"ffff0000000000000019000000000029a7fff5a700ff",
    x"ffff0000000000000001000000000029a7fff5a6f5ff",
    x"ffff0000000000000011000000000029a7fff5a6eaff",
    x"ffff0000000000000006000000000029a8fff5a6e0ff",
    x"ffff0000000000000000000000000029a7fff5a6d5ff",
    x"ffff0000000000000000000000000029a8fff5a6caff",
    x"ffff0000000000000000000000000029a8fff5a6c0ff",
    x"ffff0000000000000009000000000029a8fff5a6b5ff",
    x"ffff000000000000000a000000000029a9fff5a6aaff",
    x"ffff0000000000000011000000000029a8fff5a6a0ff",
    x"ffff000000000000001d000000000029a9fff5a695ff",
    x"ffff0000000000000012000000000029a8fff5a68aff",
    x"ffff000000000000000c000000000029a9fff5a680ff",
    x"ffff0000000000000004000000000029aafff5a675ff",
    x"ffff000000000000001d000000000029a9fff5a66aff",
    x"ffff0000000000000004000000000029a9fff5a660ff",
    x"ffff0000000000000000000000000029aafff5a655ff",
    x"ffff0000000000000000000000000029aafff5a64aff",
    x"ffff0000000000000010000000000029aafff5a63fff",
    x"ffff000000000000001e000000000029aafff5a635ff",
    x"ffff000000000000001f000000000029aafff5a62aff",
    x"ffff000000000000001f000000000029aafff5a61fff",
    x"ffff000000000000001f000000000029abfff5a615ff",
    x"ffff000000000000001f000000000029abfff5a60aff",
    x"ffff000000000000001f000000000029abfff5a5ffff",
    x"ffff000000000000001f000000000029abfff5a5f5ff",
    x"ffff000000000000001f000000000029abfff5a5eaff",
    x"ffff000000000000001f000000000029acfff5a5dfff",
    x"ffff000000000000001f000000000029abfff5a5d5ff",
    x"ffff000000000000001f000000000029acfff5a5caff",
    x"ffff000000000000001f000000000029acfff5a5bfff",
    x"ffff000000000000001f000000000029acfff5a5b5ff",
    x"ffff000000000000001f000000000029adfff5a5aaff",
    x"ffff000000000000001f000000000029acfff5a59fff",
    x"ffff000000000000001f000000000029adfff5a594ff",
    x"ffff000000000000001f000000000029adfff5a58aff",
    x"ffff000000000000001f000000000029adfff5a57fff",
    x"ffff000000000000001f000000000029adfff5a574ff",
    x"ffff000000000000001f000000000029adfff5a56aff",
    x"ffff000000000000001f000000000029aefff5a55fff",
    x"ffff000000000000001f000000000029adfff5a554ff",
    x"ffff000000000000001f000000000029aefff5a54aff",
    x"ffff000000000000001f000000000029aefff5a53fff",
    x"ffff000000000000001f000000000029aefff5a534ff",
    x"ffff000000000000001f000000000029affff5a52aff",
    x"ffff000000000000001f000000000029aefff5a51fff",
    x"ffff000000000000001f000000000029affff5a514ff",
    x"ffff000000000000001f000000000029affff5a509ff",
    x"ffff000000000000001f000000000029affff5a4ffff",
    x"ffff000000000000001f000000000029affff5a4f4ff",
    x"ffff000000000000001f000000000029affff5a4e9ff",
    x"ffff000000000000001f000000000029b0fff5a4dfff",
    x"ffff000000000000001f000000000029affff5a4d4ff",
    x"ffff000000000000001f000000000029b0fff5a4c9ff",
    x"ffff000000000000001f000000000029b0fff5a4bfff",
    x"ffff000000000000001f000000000029b0fff5a4b4ff",
    x"ffff000000000000001f000000000029b1fff5a4a9ff",
    x"ffff000000000000001f000000000029b0fff5a49fff",
    x"ffff000000000000001f000000000029b1fff5a494ff",
    x"ffff000000000000001f000000000029b1fff5a489ff",
    x"ffff0000000000000017000000000029b1fff5a47eff",
    x"ffff0000000000000006000000000029b1fff5a474ff",
    x"ffff0000000000000011000000000029b1fff5a469ff",
    x"ffff0000000000000006000000000029b2fff5a45eff",
    x"ffff0000000000000000000000000029b1fff5a454ff",
    x"ffff0000000000000000000000000029b2fff5a449ff",
    x"ffff0000000000000000000000000029b2fff5a43eff",
    x"ffff0000000000000009000000000029b3fff5a434ff",
    x"ffff000000000000000a000000000029b2fff5a429ff",
    x"ffff0000000000000011000000000029b2fff5a41eff",
    x"ffff000000000000001d000000000029b3fff5a414ff",
    x"ffff0000000000000011000000000029b3fff5a409ff",
    x"ffff0000000000000016000000000029b3fff5a3feff",
    x"ffff0000000000000005000000000029b3fff5a3f3ff",
    x"ffff0000000000000012000000000029b4fff5a3e9ff",
    x"ffff0000000000000010000000000029b3fff5a3deff",
    x"ffff0000000000000004000000000029b4fff5a3d3ff",
    x"ffff0000000000000005000000000029b4fff5a3c9ff",
    x"ffff000000000000000c000000000029b4fff5a3beff",
    x"ffff000000000000001e000000000029b4fff5a3b3ff",
    x"ffff000000000000001f000000000029b4fff5a3a9ff",
    x"ffff000000000000001b000000000029b5fff5a39eff",
    x"ffff0000000000000009000000000029b5fff5a393ff",
    x"ffff0000000000000002000000000029b5fff5a389ff",
    x"ffff000000000000001e000000000029b5fff5a37eff",
    x"ffff000000000000001d000000000029b5fff5a373ff",
    x"ffff0000000000000010000000000029b5fff5a369ff",
    x"ffff0000000000000004000000000029b6fff5a35eff",
    x"ffff0000000000000006000000000029b5fff5a353ff",
    x"ffff000000000000001f000000000029b6fff5a348ff",
    x"ffff000000000000000f000000000029b6fff5a33eff",
    x"ffff000000000000001f000000000029b7fff5a333ff",
    x"ffff000000000000001a000000000029b6fff5a328ff",
    x"ffff000000000000001b000000000029b7fff5a31eff",
    x"ffff0000000000000003000000000029b6fff5a313ff",
    x"ffff000000000000001b000000000029b7fff5a308ff",
    x"ffff000000000000000f000000000029b7fff5a2feff",
    x"ffff0000000000000016000000000029b8fff5a2f3ff",
    x"ffff000000000000001f000000000029b7fff5a2e8ff",
    x"ffff000000000000000a000000000029b8fff5a2deff",
    x"ffff000000000000001a000000000029b7fff5a2d3ff",
    x"ffff0000000000000019000000000029b8fff5a2c8ff",
    x"ffff000000000000000f000000000029b8fff5a2bdff",
    x"ffff000000000000001d000000000029b9fff5a2b3ff",
    x"ffff000000000000001b000000000029b8fff5a2a8ff",
    x"ffff0000000000000011000000000029b9fff5a29dff",
    x"ffff0000000000000003000000000029b8fff5a293ff",
    x"ffff000000000000001a000000000029b9fff5a288ff",
    x"ffff0000000000000014000000000029b9fff5a27dff",
    x"ffff000000000000000b000000000029bafff5a273ff",
    x"ffff000000000000001e000000000029b9fff5a268ff",
    x"ffff0000000000000009000000000029bafff5a25dff",
    x"ffff0000000000000009000000000029b9fff5a253ff",
    x"ffff000000000000001c000000000029bafff5a248ff",
    x"ffff000000000000001b000000000029bafff5a23dff",
    x"ffff0000000000000018000000000029bbfff5a232ff",
    x"ffff0000000000000008000000000029bafff5a228ff",
    x"ffff0000000000000006000000000029bbfff5a21dff",
    x"ffff0000000000000000000000000029bafff5a212ff",
    x"ffff0000000000000000000000000029bbfff5a208ff",
    x"ffff0000000000000018000000000029bbfff5a1fdff",
    x"ffff0000000000000004000000000029bcfff5a1f2ff",
    x"ffff0000000000000011000000000029befff5a1e8ff",
    x"ffff0000000000000006000000000029bcfff5a1ddff",
    x"ffff0000000000000000000000000029bcfff5a1d2ff",
    x"ffff0000000000000000000000000029bcfff5a1c7ff",
    x"ffff0000000000000000000000000029bcfff5a1bdff",
    x"ffff0000000000000009000000000029bcfff5a1b2ff",
    x"ffff000000000000000a000000000029bcfff5a1a7ff",
    x"ffff0000000000000011000000000029bdfff5a19dff",
    x"ffff000000000000001d000000000029bdfff5a192ff",
    x"ffff0000000000000003000000000029bdfff5a187ff"
  );
end package;